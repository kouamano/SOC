3 6
3 2 4
4 3 6
11 10 9
10 9 8
8 9 10
1 5 8
