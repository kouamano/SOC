3 4
3 2 1
4 5 6
10 9 8
1 5 8
