3 6
1 5 20
3 2 1
4 3 1
11 10 9
10 9 8
8 9 10
