5 10
A 2 3 4 5 6
B 12 13 14 5 6
C 12 13 14 15 16
D 1 1 14 5 6
E 4 1 18 7 6
F 1 3 2 5 7
G 8 17 14 15 9
H 5 1 2 5 7
I 12 10 14 7 6
J 3 2 15 7 6
