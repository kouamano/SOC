64   2000
0.964152236025835   0.3483635416653267   0.945387358826106   0.02385030656821705   0.9843629633427824   0.14273924350942932   0.1613989695592285   0.29331710461584215   0.25076792131097153   0.3453949451140481   0.3065267365692395   0.2873353913771538   0.2438111764998183   0.2667724640238826   0.30449079562757186   0.45696795315479055   0.7528680866560835   0.43539098835794   0.2048817536084007   0.27988447254786536   0.6080357275430546   0.5741286792017458   0.2410370911711503   0.3207931489903225   0.6438834915172197   0.22576513753641908   0.2956497323450443   0.29694284242210545   0.6595205281744372   0.08302589402698976   0.1342507627858158   0.0036257378062632684   0.40875260686346565   0.7376309489129417   0.8277240262165763   0.7162903464291095   0.16494143036364736   0.47085848488905907   0.5232332305890044   0.2593223932743189   0.4120733437075639   0.03546749653111904   0.3183514769806037   0.9794379207264535   0.8040376161645093   0.46133881732937326   0.07731438580945336   0.658644771736131   0.16015412464728962   0.23557367979295418   0.781664653464409   0.3617019293140256   0.5006335964728524   0.15254778576596442   0.6474138906785932   0.3580761915077623   0.09188098960938676   0.4149168368530228   0.819689864462017   0.6417858450786529   0.9269395592457395   0.9440583519639637   0.29645663387301263   0.382463451804334
0.5148662155381755   0.9085908554328447   0.978105156892409   0.4030255310778805   0.7108285993736663   0.4472520381034714   0.9007907710829556   0.7443807593417494   0.5506744747263767   0.21167835831051726   0.11912611761854654   0.3826788300277238   0.05004087825352421   0.05913057254455284   0.4717122269399533   0.024602638519961476   0.9581598886441375   0.6442137356915301   0.6520223624779363   0.3828167934413086   0.03122032939839805   0.7001553837275664   0.3555657286049237   0.00035334163697458404   0.5163541138602226   0.7915645282947217   0.37746057171251474   0.5973278105590941   0.8055255144865563   0.34431249019125026   0.47666980062955916   0.8529470512173447   0.25485103976017964   0.132634131880733   0.3575436830110126   0.4702682211896209   0.20481016150665546   0.07350355933618016   0.8858314560710593   0.44566558266965944   0.246650272862518   0.4292898236446501   0.23380909359312305   0.06284878922835084   0.21542994346411995   0.7291344399170837   0.8782433649881993   0.062495447591376256   0.6990758296038975   0.937569911622362   0.5007827932756846   0.46516763703228214   0.8935503151173412   0.5932574214311118   0.024112992646125514   0.6122205858149374   0.6386992753571614   0.4606232895503788   0.666569309635113   0.14195236462531652   0.433889113850506   0.38711973021419865   0.7807378535640536   0.6962867819556571
0.18723884098798801   0.9578299065695486   0.5469287599709306   0.6334379927273063   0.971808897523868   0.2286954666524648   0.6686853949827312   0.57094254513593   0.27273306791997065   0.29112555503010273   0.16790260170704654   0.10577490810364788   0.3791827528026295   0.6978681335989909   0.14378960906092103   0.49355432228871043   0.740483477445468   0.23724484404861212   0.4772202994258081   0.3516019576633939   0.306594363594962   0.8501251138344135   0.6964824458617546   0.6553151757077368   0.119355522606974   0.892295207264865   0.14955368589082396   0.021877182980430565   0.14754662508310595   0.6635997406124001   0.48086829090809274   0.45093463784450055   0.8748135571631354   0.37247418558229745   0.3129656892010462   0.3451597297408527   0.49563080436050583   0.6746060519833065   0.1691760801401252   0.8516054074521422   0.7551473269150378   0.4373612079346944   0.6919557807143171   0.5000034497887482   0.44855296332007577   0.5872360941002809   0.9954733348525626   0.8446882740810114   0.32919744071310175   0.694940886835416   0.8459196489617387   0.8228110911005809   0.18165081562999583   0.03134114622301578   0.36505135805364586   0.3718764532560803   0.3068372584668605   0.6588669606407184   0.05208566885259963   0.026716723515227657   0.8112064541063546   0.9842609086574118   0.8829095887124744   0.17511131606308544
0.05605912719131686   0.5468997007227174   0.19095380799815734   0.6751078662743372   0.6075061638712411   0.9596636066224365   0.19548047314559475   0.8304195921933257   0.2783087231581393   0.2647227197870206   0.34956082418385614   0.00760850109274487   0.09665790752814347   0.23338157356400482   0.9845094661302103   0.6357320478366646   0.789820649061283   0.5745146129232864   0.9324237972776107   0.6090153243214369   0.9786141949549283   0.5902537042658746   0.04951420856513623   0.43390400825835146   0.9225550677636115   0.043354003543157195   0.8585604005669789   0.7587961419840142   0.3150489038923704   0.08369039692072067   0.6630799274213841   0.9283765497906885   0.03674018073423111   0.8189676771337001   0.313519103237528   0.9207680486979436   0.9400822732060876   0.5855861035696952   0.32900963710731773   0.2850360008612791   0.15026162414480462   0.011071490646408786   0.3965858398297071   0.6760206765398422   0.1716474291898763   0.42081778638053413   0.34707163126457086   0.24211666828149075   0.2490923614262648   0.37746378283737697   0.48851123069759195   0.4833205262974765   0.9340434575338944   0.2937733859166563   0.8254313032762078   0.554943976506788   0.8973032767996633   0.47480570878295625   0.5119122000386798   0.6341759278088444   0.9572210035935756   0.8892196052132609   0.1829025629313621   0.34913992694756524
0.806959379448771   0.8781481145668522   0.786316723101655   0.673119250407723   0.6353119502588948   0.457330328186318   0.4392450918370842   0.43100258212623227   0.3862195888326299   0.07986654534894108   0.9507338611394923   0.9476820558287558   0.4521761312987355   0.7860931594322847   0.12530255786328445   0.3927380793219678   0.5548728544990722   0.31128745064932856   0.6133903578246047   0.7585621515131235   0.5976518509054966   0.4220678454360676   0.43048779489324257   0.40942222456555816   0.7906924714567255   0.5439197308692154   0.6441710717915875   0.7363029741578351   0.15538052119783075   0.08658940268289739   0.20492597995450335   0.30530039203160286   0.7691609323652008   0.006722857333956295   0.2541921188150111   0.35761833620284705   0.3169848010664653   0.2206296979016715   0.1288895609517266   0.9648802568808793   0.7621119465673931   0.9093422472523429   0.5154992031271219   0.20631810536775588   0.16446009566189657   0.48727440181627535   0.08501140823387937   0.7968958808021978   0.37376762420517107   0.9433546709470599   0.4408403364422918   0.06059290664436257   0.21838710300734035   0.8567652682641625   0.2359143564877885   0.7552925146127597   0.44922617064213954   0.8500424109302063   0.9817222376727774   0.39767417840991265   0.13224136957567423   0.6294127130285347   0.8528326767210508   0.43279392152903334
0.3701294230082811   0.7200704657761918   0.33733347359392885   0.22647581616127746   0.20566932734638457   0.23279606395991648   0.2523220653600495   0.4295799353590798   0.8319017031412135   0.2894413930128566   0.8114817289177576   0.36898702871471717   0.6135146001338732   0.43267612474869405   0.5755673724299691   0.6136945141019574   0.16428842949173364   0.5826337138184878   0.5938451347571917   0.21602033569204482   0.032047059916059405   0.9532210007899531   0.7410124580361409   0.7832264141630115   0.6619176369077783   0.23315053501376132   0.4036789844422121   0.556750598001734   0.45624830956139373   0.00035447105384482864   0.15135691908216262   0.12717066264265425   0.6243466064201803   0.7109130780409882   0.339875190164405   0.7581836339279371   0.010832006286307058   0.2782369532922942   0.7643078177344358   0.1444891198259796   0.8465435767945735   0.6956032394738064   0.17046268297724407   0.9284687841339347   0.814496516878514   0.7423822386838532   0.42945022494110313   0.1452423699709233   0.15257887997073574   0.509231703670092   0.025771240498891023   0.5884917719691892   0.6963305704093421   0.5088772326162472   0.8744143214167284   0.46132110932653503   0.07198396398916183   0.7979641545752589   0.5345391312523234   0.7031374753985979   0.06115195770285478   0.5197272012829647   0.7702313135178877   0.5586483555726184
0.21460838090828135   0.8241239618091583   0.5997686305406436   0.6301795714386835   0.40011186402976734   0.08174172312530503   0.1703184055995404   0.48493720146776026   0.24753298405903157   0.5725100194552131   0.14454716510064938   0.896445429498571   0.5512024136496895   0.06363278683896594   0.270132843683921   0.435124320172036   0.4792184496605277   0.26566863226370707   0.7355937124315975   0.731986844773438   0.4180664919576729   0.7459414309807424   0.96536239891371   0.17333848920081968   0.20345811104939154   0.921817469171584   0.36559376837306645   0.5431589177621361   0.8033462470196242   0.840075746046279   0.19527536277352603   0.05822171629437582   0.5558132629605926   0.267565726591066   0.05072819767287663   0.1617762867958048   0.004610849310903128   0.20393293975210003   0.7805953539889556   0.7266519666237689   0.5253923996503754   0.938264307488393   0.045001641557358085   0.9946651218503307   0.10732590769270253   0.1923228765076506   0.07963924264364813   0.8213266326495111   0.903867796643311   0.27050540733606654   0.7140454742705817   0.27816771488737496   0.10052154962368674   0.4304296612897875   0.5187701114970557   0.21994599859299915   0.5447082866630941   0.1628639346987215   0.46804191382417903   0.05816971179719435   0.540097437352191   0.9589309949466215   0.6874465598352234   0.3315177451734255
0.014705037701815525   0.020666687458228503   0.6424449182778653   0.33685262332309474   0.907379130009113   0.828343810950578   0.5628056756342172   0.5155259906735836   0.0035113333658020164   0.5578384036145114   0.8487602013636355   0.2373582757862087   0.9029897837421152   0.12740874232472393   0.3299900898665798   0.017412277193209515   0.3582814970790212   0.9645448076260025   0.8619481760424007   0.9592425653960152   0.8181840597268302   0.005613812679380956   0.17450161620717736   0.6277248202225897   0.8034790220250146   0.9849471252211525   0.5320566979293121   0.2908721968994949   0.8960998920159017   0.15660331427057453   0.9692510222950949   0.7753462062259112   0.8925885586500997   0.5987649106560631   0.12049082093145937   0.5379879304397025   0.9895987749079844   0.4713561683313392   0.7905007310648796   0.520575653246493   0.6313172778289632   0.5068113607053367   0.9285525550224788   0.5613330878504779   0.813133218102133   0.5011975480259558   0.7540509388153015   0.9336082676278882   0.009654196077118331   0.5162504228048034   0.2219942408859894   0.6427360707283933   0.11355430406121664   0.3596471085342288   0.25274321859089455   0.8673898645024821   0.22096574541111696   0.7608821978781657   0.1322523976594352   0.3294019340627796   0.23136697050313254   0.2895260295468265   0.34175166659455564   0.8088262808162866
0.6000496926741693   0.7827146688414898   0.41319911157207684   0.24749319296580874   0.7869164745720363   0.2815171208155339   0.6591481727567754   0.3138849253379205   0.7772622784949179   0.7652666980107306   0.43715393187078594   0.6711488546095271   0.6637079744337013   0.40561958947650173   0.1844107132798914   0.803758990107045   0.44274222902258437   0.6447373915983361   0.052158315620456204   0.4743570560442654   0.21137525851945183   0.35521136205150955   0.7104066490259006   0.6655307752279789   0.6113255658452825   0.5724966932100198   0.2972075374538238   0.41803758226217014   0.8244090912732462   0.2909795723944859   0.6380593646970484   0.10415265692424962   0.04714681277832824   0.5257128743837554   0.20090543282626247   0.43300380231472246   0.3834388383446269   0.12009328490725363   0.016494719546371068   0.6292448122076775   0.9406966093220426   0.4753558933089176   0.9643364039259149   0.154887756163412   0.7293213508025908   0.12014453125740804   0.2539297549000143   0.4893569809354332   0.11799578495730821   0.5476478380473883   0.9567222174461905   0.07131939867326302   0.293586693684062   0.2566682656529023   0.3186628527491421   0.9671667417490134   0.24643988090573377   0.730955391269147   0.11775741992287965   0.5341629394342909   0.8630010425611069   0.6108621063618933   0.10126270037650857   0.9049181272266135
0.9223044332390643   0.13550621305297575   0.1369262964505937   0.7500303710632015   0.19298308243647358   0.015361681795567714   0.8829965415505794   0.26067339012776836   0.07498729747916537   0.4677138437481795   0.9262743241043889   0.18935399145450532   0.7814006037951033   0.2110455780952772   0.6076114713552468   0.22218724970549192   0.5349607228893696   0.48009018682613025   0.48985405143236715   0.6880243102712009   0.6719596803282627   0.8692280804642369   0.38859135105585857   0.7831061830445875   0.7496552470891984   0.7337218674112612   0.2516650546052649   0.03307581198138596   0.5566721646527248   0.7183601856156935   0.36866851305468545   0.7724024218536176   0.48168486717355946   0.25064634186751394   0.44239418895029653   0.5830484303991122   0.7002842633784561   0.03960076377223676   0.8347827175950497   0.3608611806936204   0.1653235404890865   0.5595105769461065   0.3449286661626826   0.6728368704224194   0.49336386016082373   0.6902824964818696   0.956337315106824   0.8897306873778319   0.7437086130716253   0.9565606290706085   0.7046722605015591   0.856654875396446   0.1870364484189005   0.23820044345491495   0.3360037474468736   0.08425245354282836   0.705351581245341   0.987554101587401   0.8936095584965771   0.501204023143716   0.005067317866884917   0.9479533378151642   0.05882684090152737   0.1403428424500957
0.8397437773777984   0.3884427608690577   0.7138981747388448   0.4675059720276763   0.34637991721697464   0.6981602643871881   0.7575608596320208   0.5777752846498444   0.6026713041453493   0.7415996353165797   0.05288859913046176   0.7211204092533984   0.41563485572644887   0.5033991918616648   0.7168848516835882   0.6368679557105701   0.7102832744811078   0.5158450902742638   0.823275293187011   0.13566393256685397   0.7052159566142229   0.5678917524590996   0.7644484522854836   0.9953210901167583   0.8654721792364245   0.17944899159004185   0.05055027754663885   0.527815118089082   0.5190922620194498   0.4812887272028537   0.292989417914618   0.9500398334392376   0.9164209578741005   0.739689091886274   0.24010081878415623   0.2289194241858392   0.5007861021476516   0.2362899000246092   0.5232159671005682   0.5920514684752691   0.7905028276665438   0.7204448097503454   0.6999406739135571   0.4563875359084152   0.0852868710523209   0.15255305729124585   0.9354922216280734   0.4610664457916569   0.21981469181589638   0.973104065701204   0.8849419440814346   0.9332513277025749   0.7007224297964465   0.4918153384983503   0.5919525261668166   0.9832114942633374   0.784301471922346   0.7521262466120763   0.3518517073826603   0.7542920700774982   0.2835153697746944   0.5158363465874671   0.8286357402820922   0.16224060160222903
0.4930125421081506   0.7953915368371217   0.12869506636853512   0.7058530656938139   0.4077256710558297   0.6428384795458758   0.1932028447404617   0.24478661990215694   0.18791097923993327   0.6697344138446718   0.3082609006590271   0.311535292199582   0.4871885494434867   0.17791907534632154   0.7163083744922105   0.3283237979362446   0.7028870775211407   0.42579282873424523   0.3644566671095502   0.5740317278587465   0.41937170774644633   0.9099564821467782   0.5358209268274581   0.41179112625651737   0.9263591656382958   0.11456494530965647   0.4071258604589229   0.7059380605627035   0.5186334945824661   0.47172646576378063   0.21392301571846123   0.4611514406605466   0.3307225153425328   0.8019920519191088   0.9056621150594341   0.14961614846096463   0.8435339658990461   0.6240729765727873   0.18935374056722357   0.82129235052472   0.14064688837790534   0.19828014783854203   0.8248970734576733   0.24726062266597362   0.721275180631459   0.2883236656917639   0.28907614663021525   0.8354694964094562   0.7949160149931633   0.1737587203821074   0.8819502861712923   0.12953143584675272   0.27628252041069723   0.7020322546183267   0.6680272704528312   0.6683799951862062   0.9455600050681645   0.900040202699218   0.762365155393397   0.5187638467252416   0.10202603916911841   0.2759672261264307   0.5730114148261735   0.6974714962005215
0.961379150791213   0.07768707828788869   0.7481143413685002   0.45021087353454786   0.24010397015975404   0.7893634125961247   0.4590381947382849   0.6147413771250916   0.44518795516659077   0.6156046922140174   0.5770879085669925   0.4852099412783389   0.1689054347558935   0.9135724375956906   0.9090606381141614   0.8168299460921328   0.22334542968772905   0.013532234896472617   0.14669548272076438   0.2980660993668912   0.12131939051861063   0.7375650087700419   0.5736840678945909   0.6005946031663697   0.15994023972739754   0.6598779304821533   0.8255697265260908   0.15038372963182187   0.9198362695676435   0.8705145178860284   0.3665315317878059   0.5356423525067302   0.47464831440105276   0.25490982567201104   0.7894436232208134   0.05043241122839136   0.3057428796451593   0.3413373880763204   0.880382985106652   0.2336024651362586   0.08239744995743022   0.3278051531798478   0.7336875023858876   0.9355363657693674   0.9610780594388196   0.5902401444098059   0.1600034344912967   0.33494176260299763   0.8011378197114221   0.9303622139276527   0.3344337079652059   0.18455803297117576   0.8813015501437785   0.059847696041624286   0.9679021761773999   0.6489156804644455   0.40665323574272577   0.8049378703696133   0.17845855295658655   0.5984832692360541   0.1009103560975665   0.4636004822932928   0.29807556784993455   0.36488080409979556
0.018512906140136277   0.135795329113445   0.564388065464047   0.4293444383304282   0.05743484670131668   0.5455551847036391   0.40438463097275024   0.09440267572743055   0.25629702698989465   0.6151929707759863   0.06995092300754435   0.9098446427562548   0.3749954768461161   0.5553452747343621   0.1020487468301444   0.2609289622918093   0.9683422411033903   0.7504074043647488   0.9235901938735578   0.6624456930557552   0.8674318850058238   0.286806922071456   0.6255146260236233   0.2975648889559596   0.8489189788656876   0.15101159295801103   0.06112656055957635   0.8682204506255314   0.7914841321643709   0.605456408254372   0.6567419295868261   0.7738177748981009   0.5351871051744762   0.9902634374783855   0.5867910065792817   0.863973132141846   0.16019162832836015   0.43491816274402345   0.48474225974913737   0.6030441698500367   0.1918493872249698   0.6845107583792747   0.5611520658755795   0.9405984767942817   0.32441750221914595   0.3977038363078186   0.9356374398519562   0.643033587838322   0.47549852335345844   0.24669224334980758   0.8745108792923799   0.7748131372127905   0.6840143911890876   0.6412358350954356   0.2177689497055538   0.0009953623146897164   0.14882728601461132   0.6509723976170501   0.6309779431262721   0.13702223017284365   0.9886356576862512   0.2160542348730266   0.1462356833771347   0.5339780603228069
0.7967862704612814   0.531543476493752   0.5850836175015551   0.5933795835285253   0.47236876824213536   0.1338396401859334   0.6494461776495989   0.9503459956902033   0.9968702448886769   0.8871473968361258   0.774935298357219   0.17553285847741268   0.3128558536995894   0.24591156174069018   0.5571663486516653   0.17453749616272296   0.16402856768497812   0.5949391641236401   0.9261884055253932   0.03751526598987931   0.17539290999872695   0.3788849292506135   0.7799527221482585   0.5035372056670724   0.3786066395374456   0.8473414527568616   0.19486910464670332   0.9101576221385471   0.9062378712953102   0.7135018125709282   0.5454229269971044   0.9598116264483438   0.9093676264066333   0.8263544157348024   0.7704876286398854   0.7842787679709312   0.5965117727070438   0.5804428539941122   0.2133212799882202   0.6097412718082083   0.4324832050220657   0.9855036898704721   0.28713287446282704   0.5722260058183289   0.2570902950233388   0.6066187606198585   0.5071801523145686   0.06868880015125652   0.8784836554858931   0.759277307862997   0.31231104766786527   0.15853117801270936   0.9722457841905829   0.0457754952920688   0.7668881206707608   0.19871955156436547   0.06287815778394969   0.21942107955726645   0.9964004920308754   0.4144407835934343   0.4663663850769058   0.6389782255631543   0.7830792120426552   0.804699511785226
0.03388318005484009   0.6534745356926822   0.4959463375798282   0.23247350596689706   0.7767928850315013   0.04685577507282368   0.9887661852652596   0.16378470581564056   0.8983092295456081   0.2875784672098267   0.6764551375973944   0.005253527802931184   0.9260634453550252   0.2418029719177579   0.9095670169266336   0.8065339762385657   0.8631852875710755   0.022381892360491474   0.9131665248957581   0.3920931926451314   0.3968189024941697   0.38340366679733723   0.1300873128531029   0.5873936808599054   0.3629357224393296   0.729929131104655   0.6341409752732747   0.35492017489300837   0.5861428374078282   0.6830733560318313   0.6453747900080151   0.1911354690773678   0.6878336078622201   0.3954948888220046   0.9689196524106207   0.1858819412744366   0.761770162507195   0.15369191690424672   0.05935263548398716   0.3793479650358709   0.8985848749361195   0.13131002454375526   0.14618611058822903   0.9872547723907394   0.5017659724419499   0.747906357746418   0.01609879773512615   0.39986109153083405   0.13883025000262028   0.01797722664176302   0.38195782246185145   0.04494091663782569   0.552687412594792   0.3349038706099317   0.7365830324538364   0.8538054475604578   0.8648538047325719   0.9394089817879271   0.7676633800432157   0.6679235062860213   0.10308364222537687   0.7857170648836803   0.7083107445592285   0.28857554125015034
0.20449876728925737   0.6544070403399251   0.5621246339709994   0.3013207688594109   0.7027327948473076   0.906500682593507   0.5460258362358733   0.9014596773285768   0.5639025448446873   0.8885234559517441   0.16406801377402186   0.8565187606907512   0.011215132249895244   0.5536195853418123   0.42748498132018553   0.0027133131302932564   0.1463613275173234   0.6142106035538853   0.6598216012769699   0.334789806844272   0.04327768529194651   0.8284935386702049   0.9515108567177414   0.04621426559412163   0.8387789180026891   0.17408649833027987   0.3893862227467419   0.7448934967347107   0.13604612315538162   0.2675858157367728   0.8433603865108686   0.8434338194061339   0.5721435783106944   0.3790623597850288   0.6792923727368467   0.9869150587153828   0.5609284460607992   0.8254427744432165   0.2518073914166612   0.9842017455850895   0.4145671185434757   0.21123217088933113   0.5919857901396913   0.6494119387408175   0.3712894332515292   0.3827386322191262   0.64047493342195   0.6031976731466959   0.5325105152488401   0.2086521338888463   0.2510887106752081   0.8583041764119852   0.39646439209345846   0.9410663181520734   0.4077283241643395   0.014870357005851233   0.8243208137827641   0.5620039583670446   0.7284359514274928   0.02795529829046847   0.263392367721965   0.7365611839238283   0.4766285600108316   0.04375355270537896
0.8488252491784892   0.5253290130344971   0.8846427698711402   0.3943416139645614   0.47753581592696004   0.14259038081537093   0.2441678364491902   0.7911439408178655   0.94502530067812   0.9339382469265246   0.993079125773982   0.9328397644058805   0.5485609085846616   0.9928719287744512   0.5853508016096426   0.9179694074000292   0.7242400948018974   0.4308679704074065   0.8569148501821497   0.8900141091095607   0.46084772707993243   0.6943067864835782   0.38028629017131815   0.8462605564041817   0.6120224779014432   0.1689777734490811   0.4956435203001779   0.45191894243962033   0.1344866619744831   0.026387392633710174   0.2514756838509877   0.6607750016217547   0.18946136129636312   0.09244914570718554   0.2583965580770056   0.7279352372158744   0.6409004527117016   0.09957721693273439   0.6730457564673631   0.8099658298158452   0.9166603579098042   0.6687092465253279   0.8161309062852133   0.9199517207062845   0.4558126308298718   0.9744024600417497   0.43584461611389524   0.07369116430210275   0.8437901529284286   0.8054246865926686   0.9402010958137174   0.6217722218624825   0.7093034909539455   0.7790372939589584   0.6887254119627296   0.9609972202407276   0.5198421296575824   0.6865881482517728   0.430328853885724   0.23306198302485334   0.8789416769458808   0.5870109313190385   0.7572830974183609   0.4230961532090081
0.9622813190360766   0.9183016847937105   0.9411521911331475   0.5031444325027237   0.5064686882062048   0.9438992247519609   0.5053075750192523   0.4294532682006209   0.6626785352777762   0.13847453815929228   0.565106479205535   0.8076810463381384   0.9533750443238307   0.35943724420033385   0.8763810672428054   0.8466838260974108   0.43353291466624827   0.672849095948561   0.4460522133570814   0.6136218430725574   0.5545912377203674   0.08583816462952251   0.6887691159387205   0.19052568986354929   0.592309918684291   0.16753647983581194   0.7476169248055728   0.6873812573608257   0.08584123047808614   0.22363725508385107   0.24230934978632057   0.25792798916020476   0.42316269520030997   0.08516271692455878   0.6772028705807855   0.4502469428220663   0.46978765087647933   0.7257254727242249   0.8008218033379803   0.6035631167246555   0.0362547362102311   0.052876376775663904   0.35476958998089886   0.989941273652098   0.4816634984898636   0.9670382121461414   0.6660004740421784   0.7994155837885487   0.8893535798055727   0.7995017323103295   0.9183835492366055   0.11203432642772312   0.8035123493274865   0.5758644772264784   0.6760741994502849   0.8541063372675184   0.38034965412717653   0.49070176030191964   0.9988713288694994   0.4038593944454521   0.9105620032506971   0.7649762875776948   0.1980495255315191   0.8002962777207966
0.8743072670404661   0.7120999108020308   0.8432799355506203   0.8103550040686985   0.39264376855060246   0.7450616986558894   0.17727946150844187   0.01093942028014977   0.5032901887450298   0.9455599663455599   0.2588959122718364   0.8989050938524267   0.6997778394175432   0.36969548911908157   0.5828217128215515   0.04479875658490826   0.31942818529036676   0.878993728817162   0.5839503839520521   0.6409393621394561   0.40886618203966957   0.11401744123946722   0.38590085842053307   0.8406430844186595   0.5345589149992035   0.4019175304374364   0.5426209228699128   0.030288080349961027   0.14191514644860098   0.6568558317815469   0.3653414613614709   0.019348660069811258   0.6386249577035712   0.711295865435987   0.1064455490896345   0.12044356621738461   0.938847118286028   0.34160037631690543   0.523623836268083   0.07564480963247634   0.6194189329956612   0.46260664749974345   0.9396734523160308   0.4347054474930202   0.21055275095599163   0.3485892062602763   0.5537725938954978   0.5940623630743607   0.6759938359567882   0.9466716758228398   0.01115167102558504   0.5637742827243996   0.5340786895081872   0.2898158440412929   0.6458102096641142   0.5444256226545884   0.895453731804616   0.5785199786053059   0.5393646605744796   0.4239820564372037   0.9566066135185881   0.23691960228840048   0.015740824306396662   0.3483372468047274
0.3371876805229269   0.774312954788657   0.07606737199036581   0.9136317993117072   0.12663492956693528   0.42572374852838074   0.522294778094868   0.31956943623734657   0.45064109361014715   0.4790520727055409   0.511143107069283   0.755795153512947   0.91656240410196   0.189236228664248   0.8653328974051688   0.21136953085835863   0.021108672297343978   0.610716250058942   0.32596823683068915   0.7873874744211549   0.0645020587787559   0.3737966477705416   0.3102274125242925   0.43905022761642754   0.727314378255829   0.5994836929818845   0.23416004053392667   0.5254184283047203   0.6006794486888937   0.17375994445350382   0.7118652624390587   0.20584899206737375   0.15003835507874658   0.694707871747963   0.2007221553697757   0.45005383855442677   0.2334759509767866   0.505471643083715   0.3353892579646069   0.23868430769606813   0.21236727867944263   0.8947553930247729   0.009421021133917733   0.4512968332749132   0.14786521990068674   0.5209587452542312   0.6991936086096252   0.012246605658485687   0.42055084164485773   0.9214750522723467   0.46503356807569857   0.4868281773537653   0.819871392955964   0.7477151078188429   0.75316830563664   0.2809791852863916   0.6698330378772175   0.05300723607087994   0.5524461502668643   0.8309253467319648   0.43635708690043085   0.547535592987165   0.21705689230225736   0.5922410390358966
0.22398980822098824   0.6527801999623921   0.20763587116833962   0.14094420576098343   0.07612458832030151   0.13182145470816078   0.5084422625587144   0.12869760010249773   0.6555737466754438   0.21034640243581407   0.043408694483015785   0.6418694227487324   0.8357023537194798   0.46263129461697117   0.2902403888463759   0.36089023746234083   0.16586931584226225   0.40962405854609124   0.7377942385795117   0.529964890730376   0.7295122289418314   0.8620884655589263   0.5207373462772543   0.9377238516944794   0.5055224207208432   0.20930826559653418   0.3131014751089147   0.7967796459334959   0.42939783240054163   0.07748681088837338   0.8046592125502003   0.6680820458309982   0.7738240857250979   0.8671404084525594   0.7612505180671845   0.026212623082265827   0.9381217320056181   0.40450911383558813   0.47101012922080865   0.6653223856199251   0.7722524161633559   0.9948850552894969   0.733215890641297   0.135357494889549   0.0427401872215245   0.13279658973057062   0.21247854436404273   0.19763364319506962   0.5372177665006813   0.9234883241340365   0.8993770692551281   0.40085399726157367   0.10781993410013971   0.8460015132456631   0.09471785670492777   0.7327719514305755   0.3339958483750418   0.9788611047931037   0.33346733863774325   0.7065593283483096   0.3958741163694237   0.5743519909575157   0.8624572094169346   0.041236942728384615
0.6236217002060678   0.5794669356680188   0.1292413187756376   0.9058794478388356   0.5808815129845433   0.44667034593744814   0.9167627744115949   0.708245804643766   0.04366374648386197   0.5231820218034117   0.01738570515646681   0.3073918073821923   0.9358438123837223   0.6771805085577486   0.922667848451539   0.5746198559516168   0.6018479640086805   0.6983194037646447   0.5892005098137958   0.8680605276033072   0.20597384763925672   0.12396741280712914   0.7267433003968612   0.8268235848749226   0.5823521474331889   0.5445004771391104   0.5975019816212236   0.920944137036087   0.001470634448645579   0.09783013120166226   0.6807392072096287   0.212698332392321   0.9578068879647836   0.5746481093982506   0.6633535020531619   0.9053065250101286   0.021963075581061357   0.897467600840502   0.7406856536016229   0.33068666905851185   0.42011511157238096   0.19914819707585726   0.15148514378782704   0.46262614145520464   0.21414126393312424   0.07518078426872812   0.4247418433909659   0.6358025565802821   0.6317891164999353   0.5306803071296178   0.8272398617697424   0.714858419544195   0.6303184820512897   0.4328501759279555   0.14650065456011369   0.5021600871518741   0.6725115940865062   0.8582020665297049   0.48314715250695184   0.5968535621417453   0.6505485185054448   0.9607344656892028   0.742461498905329   0.2661668930832335
0.23043340693306386   0.7615862686133456   0.5909763551175019   0.8035407516280288   0.016292142999939606   0.6864054843446175   0.16623451172653606   0.16773819504774684   0.3845030265000043   0.1557251772149997   0.3389946499567937   0.4528797755035518   0.7541845444487145   0.7228750012870442   0.19249399539668   0.9507196883516777   0.08167295036220835   0.8646729347573393   0.7093468428897282   0.3538661262099324   0.4311244318567636   0.9039384690681365   0.9668853439843992   0.08769923312669888   0.20069102492369972   0.1423522004547909   0.3759089888668972   0.28415848149867   0.1843988819237601   0.45594671611017346   0.20967447714036117   0.11642028645092317   0.7998958554237559   0.3002215388951738   0.8706798271835675   0.6635405109473714   0.045711310975041344   0.5773465376081296   0.6781858317868875   0.7128208225956937   0.964038360612833   0.7126736028507903   0.9688389888971592   0.3589546963857613   0.5329139287560694   0.8087351337826537   0.00195364491276012   0.2712554632590624   0.3322229038323697   0.6663829333278628   0.6260446560458629   0.9870969817603924   0.14782402190860955   0.21043621721768938   0.41637017890550176   0.8706766953094692   0.3479281664848537   0.9102146783225156   0.5456903517219343   0.20713618436209782   0.30221685550981237   0.33286814071438603   0.8675045199350468   0.49431536176640417
0.3381784948969794   0.6201945378635958   0.8986655310378875   0.13536066538064292   0.80526456614091   0.811459404080942   0.8967118861251274   0.8641052021215805   0.4730416623085403   0.14507647075307914   0.2706672300792645   0.8770082203611882   0.32521764039993073   0.9346402535353898   0.8542970511737628   0.006331525051718936   0.977289473915077   0.02442557521287417   0.3086066994518285   0.7991953406896211   0.6750726184052647   0.6915574344984882   0.44110217951678166   0.30487997892321694   0.3368941235082853   0.0713628966348924   0.5424366484788942   0.16951931354257402   0.5316295573673753   0.2599034925539504   0.6457247623537667   0.3054141114209935   0.058587895058835035   0.11482702180087126   0.3750575322745022   0.4284058910598053   0.7333702546589043   0.1801867682654815   0.5207604811007395   0.4220743660080864   0.7560807807438272   0.15576119305260733   0.21215378164891102   0.6228790253184653   0.08100816233856262   0.46420375855411916   0.7710516021321293   0.31799904639524834   0.7441140388302774   0.3928408619192268   0.2286149536532352   0.14847973285267435   0.21248448146290203   0.13293736936527636   0.5828901912994685   0.8430656214316808   0.15389658640406698   0.018110347564405112   0.20783265902496623   0.41465973037187553   0.4205263317451627   0.8379235792989236   0.6870721779242267   0.9925853643637892
0.6644455510013354   0.6821623862463163   0.47491839627531574   0.36970633904532385   0.5834373886627727   0.21795862769219712   0.7038667941431864   0.051707292650075495   0.8393233498324955   0.8251177657729704   0.47525184048995117   0.9032275597974011   0.6268388683695935   0.692180396407694   0.8923616491904827   0.06016193836572028   0.47294228196552646   0.6740700488432889   0.6845289901655165   0.6455022079938447   0.05241595022036376   0.8361464695443652   0.9974568122412898   0.6529168436300556   0.3879703992190284   0.15398408329804897   0.5225384159659741   0.28321050458473174   0.8045330105562556   0.9360254556058518   0.8186716218227876   0.23150321193465626   0.9652096607237601   0.11090768983288148   0.3434197813328365   0.32827565213725507   0.3383707923541667   0.4187272934251875   0.4510581321423538   0.2681137137715348   0.8654285103886403   0.7446572445818986   0.7665291419768373   0.6226115057776901   0.8130125601682765   0.9085107750375334   0.7690723297355475   0.9696946621476344   0.4250421609492482   0.7545266917394844   0.24653391376957348   0.6864841575629027   0.6205091503929926   0.8185012361336326   0.4278622919467858   0.4549809456282465   0.6552994896692325   0.7075935463007511   0.08444251061394932   0.1267052934909914   0.31692869731506573   0.28886625287556356   0.6333843784715956   0.8585915797194565
0.45150018692642546   0.5442090082936649   0.8668552364947583   0.2359800739417665   0.638487626758149   0.6356982332561316   0.09778290675921074   0.266285411794132   0.21344546580890075   0.8811715415166472   0.8512489929896373   0.5798012542312293   0.5929363154159082   0.06267030538301464   0.4233867010428514   0.12482030860298278   0.9376368257466757   0.35507675908226355   0.3389441904289021   0.9981150151119914   0.62070812843161   0.06621050620669999   0.7055598119573065   0.13952343539253478   0.1692079415051846   0.5220014979130351   0.8387045754625483   0.9035433614507683   0.5307203147470356   0.8863032646569035   0.7409216687033376   0.6372579496566363   0.3172748489381349   0.005131723140256225   0.8896726757137003   0.057456695425406996   0.7243385335222268   0.9424614177572416   0.46628597467084887   0.9326363868224242   0.7867017077755509   0.587384658674978   0.12734178424194675   0.9345213717104328   0.16599357934394096   0.521174152468278   0.4217819722846402   0.7949979363178981   0.9967856378387564   0.999172654555243   0.5830773968220918   0.8914545748671298   0.4660653230917207   0.11286938989833957   0.8421557281187543   0.25419662521049347   0.14879047415358584   0.10773766675808334   0.9524830524050539   0.19673992978508648   0.4244519406313591   0.16527624900084176   0.48619707773420506   0.26410354296266225
0.6377502328558081   0.5778915903258638   0.35885529349225825   0.32958217125222944   0.4717566535118672   0.05671743785758573   0.9370733212076181   0.5345842349343314   0.4749710156731108   0.05754478330234272   0.35399592438552624   0.6431296600672016   0.00890569258139004   0.9446753934040032   0.511840196266772   0.38893303485670816   0.8601152184278043   0.8369377266459198   0.5593571438617181   0.19219310507162166   0.4356632777964451   0.671661477645078   0.073160066127513   0.9280895621089593   0.797913044940637   0.09376988731921429   0.7143047726352547   0.59850739085673   0.3261563914287698   0.03705244946162857   0.7772314514276366   0.06392315592239857   0.851185375755659   0.9795076661592859   0.4232355270421104   0.42079349585519693   0.842279683174269   0.03483227275528269   0.9113953307753384   0.03186046099848881   0.9821644647464648   0.19789454610936288   0.3520381869136204   0.8396673559268671   0.5465011869500197   0.5262330684642849   0.2788781207861074   0.9115777938179078   0.7485881420093827   0.43246318114507054   0.5645733481508527   0.31307040296117783   0.42243175058061294   0.395410731683442   0.7873418967232161   0.24914724703877927   0.5712463748249539   0.4159030655241561   0.36410636968110566   0.8283537511835823   0.7289666916506848   0.38107079276887346   0.4527110389057672   0.7964932901850935
0.7468022269042202   0.18317624665951057   0.1006728519921468   0.9568259342582264   0.20030103995420043   0.6569431781952257   0.8217947312060394   0.04524814044031856   0.45171289794481767   0.22447999705015517   0.2572213830551867   0.7321777374791407   0.029281147364204778   0.8290692653667132   0.4698794863319707   0.48303049044036145   0.4580347725392509   0.41316619984255704   0.10577311665086506   0.6546767392567792   0.729068080888566   0.03209540707368361   0.6530620777450978   0.8581834490716856   0.9822658539843458   0.848919160414173   0.552389225752951   0.9013575148134593   0.7819648140301455   0.19197598221894732   0.7305944945469116   0.8561093743731407   0.3302519160853278   0.9674959851687921   0.4733731114917249   0.12393163689399998   0.300970768721123   0.13842671980207893   0.0034936251597542265   0.6409011464536385   0.8429359961818721   0.7252605199595219   0.8977205085088892   0.9862244071968594   0.11386791529330612   0.6931651128858383   0.24465843076379132   0.12804095812517383   0.1316020613089602   0.8442459524716652   0.6922692050108402   0.22668344331171458   0.34963724727881473   0.6522699702527179   0.9616747104639286   0.3705740689385739   0.01938533119348694   0.6847739850839258   0.4883015989722037   0.24664243204457392   0.7184145624723639   0.5463472652818469   0.48480797381244944   0.6057412855909354
0.8754785662904918   0.821086745322325   0.5870874653035603   0.619516878394076   0.7616106509971857   0.12792163243648672   0.342429034539769   0.49147592026890213   0.6300085896882255   0.28367567996482146   0.6501598295289287   0.26479247695718755   0.28037134240941075   0.6314057097121035   0.6884851190650001   0.8942184080186136   0.2609860112159238   0.9466317246281777   0.2001835200927964   0.6475759759740397   0.5425714487435599   0.4002844593463309   0.7153755462803469   0.04183469038310433   0.6670928824530681   0.5791977140240059   0.12828808097678665   0.4223178119890284   0.9054822314558824   0.4512760815875192   0.7858590464370176   0.9308418917201262   0.27547364176765693   0.16760040162269774   0.13569921690808895   0.6660494147629388   0.9951022993582462   0.5361946919105942   0.44721409784308885   0.7718310067443251   0.7341162881423224   0.5895629672824164   0.2470305777502924   0.1242550307702854   0.19154483939876255   0.18927850793608558   0.5316550314699454   0.08242034038718106   0.5244519569456945   0.6100807939120797   0.4033669504931588   0.6601025283981526   0.6189697254898121   0.15880471232456048   0.6175079040561412   0.7292606366780264   0.3434960837221552   0.9912043107018628   0.4818086871480522   0.0632112219150877   0.348393784363909   0.45500961879126856   0.03459458930496337   0.29138021517076257
0.6142774962215866   0.8654466515088521   0.7875640115546709   0.1671251844004772   0.422732656822824   0.6761681435727666   0.25590898008472546   0.08470484401329613   0.8982806998771296   0.06608734966068686   0.8525420295915667   0.42460231561514344   0.2793109743873174   0.9072826373361264   0.23503412553542552   0.6953416789371171   0.9358148906651622   0.9160783266342636   0.7532254383873733   0.6321304570220293   0.5874211063012532   0.4610687078429951   0.7186308490824099   0.34075024185126673   0.9731436100796667   0.595622056334143   0.931066837527739   0.17362505745078952   0.5504109532568426   0.9194539127613764   0.6751578574430135   0.08892021343749339   0.6521302533797131   0.8533665631006896   0.8226158278514468   0.66431789782235   0.3728192789923957   0.9460839257645632   0.5875817023160214   0.9689762188852329   0.4370043883272335   0.030005599130299564   0.834356263928648   0.3368457618632036   0.8495832820259802   0.5689368912873045   0.11572541484623806   0.9960955200119369   0.8764396719463136   0.9733148349531615   0.18465857731849908   0.8224704625611473   0.3260287186894709   0.0538609221917851   0.5095007198754856   0.733550249123654   0.6738984653097578   0.20049435909109553   0.6868848920240387   0.06923235130130402   0.3010791863173621   0.25441043332653235   0.09930318970801742   0.1002561324160711
0.8640747979901287   0.22440483419623278   0.2649469257793694   0.7634103705528675   0.014491515964148341   0.6554679429089283   0.14922151093313135   0.7673148505409306   0.13805184401783474   0.6821531079557668   0.9645629336146323   0.9448443879797833   0.8120231253283638   0.6282921857639816   0.4550622137391467   0.2112941388561293   0.13812466001860602   0.42779782667288613   0.768177321715108   0.1420617875548253   0.8370454737012439   0.17338739334635378   0.6688741320070906   0.04180565513875417   0.9729706757111153   0.948982559150121   0.40392720622772116   0.2783952845858867   0.958479159746967   0.29351461624119274   0.2547056952945898   0.5110804340449561   0.8204273157291322   0.611361508285426   0.2901427616799575   0.5662360460651727   0.008404190400768407   0.9830693225214443   0.8350805479408108   0.35494190720904345   0.8702795303821624   0.5552714958485582   0.06690322622570286   0.2128801196542182   0.033234056680918486   0.38188410250220445   0.3980290942186123   0.17107446451546401   0.060263380969803174   0.4329015433520834   0.9941018879908912   0.8926791799295773   0.1017842212228362   0.13938692711089068   0.7393961926963014   0.3815987458846213   0.28135690549370396   0.5280254188254647   0.44925343101634385   0.8153626998194485   0.27295271509293556   0.5449560963040203   0.6141728830755331   0.460420792610405
0.4026731847107732   0.9896846004554621   0.5472696568498302   0.24754067295618687   0.3694391280298547   0.6078004979532577   0.14924056263121788   0.07646620844072284   0.3091757470600515   0.17489895460117427   0.1551386746403267   0.18378702851114548   0.20739152583721532   0.035512027490283614   0.4157424819440253   0.8021882826265242   0.9260346203435114   0.507486608664819   0.9664890509276814   0.9868255828070757   0.6530819052505757   0.9625305123607986   0.3523161678521484   0.5264047901966706   0.25040872053980257   0.9728459119053365   0.8050465110023182   0.27886411724048377   0.8809695925099479   0.3650454139520788   0.6558059483711003   0.2023979087997609   0.5717938454498964   0.1901464593509045   0.5006672737307736   0.018610880288615426   0.3644023196126811   0.1546344318606209   0.0849247917867483   0.21642259766209124   0.43836769926916974   0.647147823195802   0.11843574085906684   0.22959701485501557   0.785285794018594   0.6846173108350033   0.7661195730069185   0.703192224658345   0.5348770734787914   0.7117713989296669   0.9610730620046002   0.4243281074178612   0.6539074809688435   0.34672598497758805   0.3052671136334999   0.2219301986181003   0.0821136355189471   0.15657952562668356   0.8045998399027263   0.20331931832948485   0.717711315906266   0.0019450937660626868   0.7196750481159779   0.9868967206673936
0.2793436166370962   0.3547972705702607   0.6012393072569111   0.757299705812378   0.49405782261850223   0.6701799597352573   0.8351197342499926   0.0541074811540331   0.9591807491397109   0.9584085608055906   0.8740466722453925   0.6297793737361719   0.30527326817086736   0.6116825758280025   0.5687795586118926   0.4078491751180716   0.22315963265192026   0.45510305020131886   0.7641797187091662   0.2045298567885868   0.5054483167456543   0.4531579564352562   0.044504670593188314   0.21763313612119317   0.22610470010855802   0.09836068586499545   0.4432653633362772   0.46033343030881513   0.7320468774900558   0.42818072612973807   0.6081456290862846   0.406225949154782   0.772866128350345   0.4697721653241475   0.7340989568408921   0.7764465754186101   0.46759286017947754   0.8580895894961451   0.1653193982289995   0.3685974003005385   0.2444332275275573   0.4029865392948262   0.4011396795198332   0.16406754351195169   0.7389849107819031   0.94982858285957   0.3566350089266449   0.9464344073907586   0.512880210673345   0.8514678969945746   0.9133696455903677   0.48610097708194344   0.7808333331832893   0.42328717086483647   0.3052240165040832   0.0798750279271614   0.007967204832944363   0.9535150055406889   0.5711250596631912   0.30342845250855127   0.5403743446534668   0.09542541604454388   0.40580566143419167   0.9348310522080128
0.2959411171259095   0.6924388767497177   0.004665981914358448   0.7707635086960611   0.5569562063440064   0.7426102938901477   0.6480309729877135   0.8243291013053026   0.04407599567066137   0.8911423968955732   0.7346613273973458   0.3382281242233592   0.2632426624873721   0.46785522603073665   0.42943731089326265   0.2583530962961978   0.2552754576544277   0.5143402204900477   0.8583122512300715   0.9549246437876465   0.7149011130009609   0.41891480444550383   0.4525065897958799   0.020093591579633665   0.41895999587505145   0.7264759276957862   0.4478406078815214   0.24933008288357256   0.8620037895310451   0.9838656338056385   0.7998096348938079   0.42500098157826993   0.8179277938603836   0.09272323691006532   0.065148307496462   0.08677285735491078   0.5546851313730116   0.6248680108793286   0.6357109966031993   0.828419761058713   0.29940967371858385   0.11052779038928094   0.7773987453731278   0.8734951172710665   0.5845085607176229   0.6916129859437771   0.324892155577248   0.8534015256914329   0.16554856484257147   0.9651370582479909   0.8770515476957266   0.6040714428078603   0.3035447753115264   0.9812714244423525   0.07724191280191872   0.17907046122959036   0.48561698145114274   0.8885481875322871   0.012093605305456716   0.09229760387467958   0.9309318500781312   0.2636801766529585   0.37638260870225737   0.2638778428159666
0.6315221763595473   0.15315238626367755   0.5989838633291296   0.39038272554490006   0.047013615641924425   0.4615394003199005   0.2740917077518816   0.5369811998534672   0.881465050799353   0.49640234207190953   0.397040160056155   0.9329097570456069   0.5779202754878265   0.5151309176295571   0.3197982472542363   0.7538392958160165   0.0923032940366838   0.62658273009727   0.30770464194877956   0.6615416919413369   0.16137144395855263   0.3629025534443114   0.9313220332465222   0.39766384912537034   0.5298492675990053   0.20975016718063383   0.3323381699173927   0.007281123580470298   0.4828356519570809   0.7482107668607334   0.05824646216551109   0.47029992372700313   0.6013706011577279   0.2518084247888238   0.661206302109356   0.5373901666813963   0.023450325669901344   0.7366775071592667   0.3414080548551198   0.7835508708653798   0.9311470316332175   0.11009477706199688   0.033703412906340255   0.12200917892404282   0.7697755876746649   0.7471922236176854   0.10238137965981807   0.7243453297986725   0.23992632007565962   0.5374420564370517   0.7700432097424255   0.7170642062182022   0.7570906681185787   0.7892312895763183   0.7117967475769144   0.24676428249119906   0.15572006696085086   0.5374228647874945   0.05059044546755823   0.7093741158098028   0.1322697412909495   0.8007453576282277   0.7091823906124384   0.925823244944423
0.20112270965773196   0.6906505805662309   0.6754789777060981   0.8038140660203803   0.43134712198306707   0.9434583569485453   0.5730975980462801   0.07946873622170778   0.19142080190740743   0.4060163005114937   0.8030543883038547   0.3624045300035056   0.4343301337888287   0.6167850109351753   0.09125764072694034   0.11564024751230653   0.27861006682797784   0.07936214614768089   0.040667195259382116   0.4062661317025037   0.1463403255370283   0.2786167885194532   0.3314848046469437   0.48044288675808067   0.9452176158792963   0.5879662079532224   0.6560058269408455   0.6766288207377004   0.5138704938962293   0.644507851004677   0.08290822889456546   0.5971600845159926   0.32244969198882184   0.23849155049318335   0.2798538405907108   0.234755554512487   0.8881195581999931   0.6217065395580079   0.18859619986377044   0.11911530700018047   0.6095094913720154   0.542344393410327   0.14792900460438832   0.7128491752976768   0.463169165834987   0.2637276048908739   0.8164441999574447   0.2324062885395961   0.5179515499556907   0.6757613969376515   0.16043837301659908   0.5557774678018957   0.004081056059461454   0.03125354593297449   0.0775301441220336   0.9586173832859031   0.6816313640706396   0.7927619954397912   0.7976763035313228   0.7238618287734161   0.7935118058706465   0.17105545588178317   0.6090801036675524   0.6047465217732356
0.18400231449863114   0.6287110624714561   0.4611510990631641   0.8918973464755588   0.7208331486636441   0.3649834575805822   0.6447068991057194   0.6594910579359627   0.20288159870795336   0.6892220606429307   0.4842685260891204   0.10371359013406706   0.1988005426484919   0.6579685147099562   0.4067383819670868   0.14509620684816396   0.5171691785778523   0.8652065192701651   0.609062078435764   0.42123437807474784   0.7236573727072059   0.6941510633883818   0.9999819747682116   0.8164878563015122   0.5396550582085747   0.06544000091692578   0.5388308757050475   0.9245905098259533   0.8188219095449306   0.7004565433363436   0.8941239765993281   0.2650994518899905   0.6159403108369772   0.011234482693412862   0.40985545051020766   0.16138586175592345   0.41713976818848536   0.35326596798345666   0.003117068543120876   0.016289654907759507   0.899970589610633   0.4880594487132916   0.3940549901073569   0.5950552768330116   0.17631321690342724   0.7939083853249097   0.39407301533914535   0.7785674205314995   0.6366581586948525   0.7284683844079839   0.8552421396340979   0.8539769107055462   0.8178362491499219   0.02801184107164034   0.9611181630347698   0.5888774588155556   0.2018959383129447   0.016777358378227476   0.5512627125245622   0.4274915970596322   0.7847561701244593   0.6635113903947708   0.5481456439814413   0.41120194215187267
0.8847855805138263   0.17545194168147923   0.15409065387408435   0.816146665318861   0.708472363610399   0.38154355635656956   0.760017638534939   0.03757924478736155   0.07181420491554646   0.6530751719485857   0.9047754989008412   0.18360233408181537   0.25397795576562454   0.6250633308769453   0.9436573358660714   0.5947248752662597   0.05208201745267983   0.6082859724987179   0.3923946233415092   0.16723327820662753   0.2673258473282205   0.944774582103947   0.8442489793600679   0.7560313360547548   0.38254026681439424   0.7693226404224678   0.6901583254859837   0.9398846707358938   0.6740679032039952   0.3877790840658982   0.9301406869510446   0.9023054259485322   0.6022536982884488   0.7347039121173126   0.025365188050203463   0.7187030918667169   0.3482757425228242   0.10964058124036725   0.08170785218413211   0.12397821660045717   0.2961937250701444   0.5013546087416494   0.6893132288426229   0.9567449383938297   0.028867877741923904   0.5565800266377025   0.8450642494825549   0.20071360233907481   0.6463276109275297   0.7872573862152347   0.1549059239965713   0.260828931603181   0.9722597077235344   0.39947830214933644   0.2247652370455267   0.35852350565464874   0.3700060094350857   0.6647743900320239   0.19940004899532324   0.6398204137879319   0.021730266912261452   0.5551338087916566   0.11769219681119113   0.5158421971874747
0.725536541842117   0.0537792000500072   0.4283789679685682   0.559097258793645   0.6966686641001931   0.4971991734123048   0.5833147184860134   0.3583836564545702   0.05034105317266348   0.7099417871970701   0.428408794489442   0.0975547248513892   0.07808134544912902   0.3104634850477337   0.20364355744391532   0.7390312191967404   0.7080753360140434   0.6456890950157098   0.004243508448592084   0.09921080540880861   0.6863450691017818   0.0905552862240532   0.886551311637401   0.583368608221334   0.9608085272596648   0.036776086174046   0.4581723436688327   0.02427134942768889   0.2641398631594717   0.5395769127617412   0.8748576251828194   0.6658876929731187   0.2137988099868082   0.8296351255646711   0.4464488306933774   0.5683329681217295   0.1357174645376792   0.5191716405169374   0.24280527324946208   0.829301748924989   0.42764212852363587   0.8734825455012275   0.23856176480087   0.7300909435161804   0.741297059421854   0.7829272592771743   0.352010453163469   0.14672233529484646   0.7804885321621892   0.7461511731031284   0.8938381094946363   0.12245098586715758   0.5163486690027175   0.20657426034138712   0.01898048431181692   0.4565632928940389   0.30254985901590925   0.37693913477671603   0.5725316536184395   0.8882303247723095   0.16683239447823006   0.8577674942597787   0.32972638036897745   0.05892857584732043
0.7391902659545942   0.9842849487585511   0.09116461556810743   0.32883763233114005   0.9978932065327403   0.20135768948137678   0.7391541624046384   0.18211529703629356   0.2174046743705511   0.45520651637824844   0.8453160529100021   0.05966431116913598   0.7010560053678336   0.24863225603686132   0.8263355685981851   0.6031010182750971   0.3985061463519244   0.8716931212601452   0.25380391497974564   0.7148706935027876   0.23167375187369432   0.013925627000366564   0.9240775346107682   0.6559421176554672   0.49248348591910013   0.02964067824181543   0.8329129190426607   0.3271044853243272   0.49459027938635985   0.8282829887604386   0.09375875663802238   0.14498918828803362   0.27718560501580874   0.3730764723821902   0.24844270372802033   0.08532487711889762   0.576129599647975   0.12444421634532889   0.42210713512983516   0.48222385884380053   0.1776234532960507   0.2527510950851836   0.16830322015008953   0.7673531653410129   0.9459497014223563   0.23882546808481708   0.24422568553932134   0.1114110476855457   0.4534662155032563   0.20918478984300165   0.4113127664966606   0.7843065623612185   0.9588759361168964   0.380901801082563   0.3175540098586382   0.6393173740731849   0.6816903311010877   0.00782532870037281   0.06911130613061787   0.5539924969542873   0.10556073145311254   0.8833811123550439   0.6470041710007827   0.07176863811048675
0.9279372781570618   0.6306300172698603   0.47870095085069314   0.30441547276947384   0.9819875767347055   0.3918045491850432   0.2344752653113718   0.19300442508392815   0.5285213612314492   0.18261975934204158   0.8231624988147113   0.40869786272270964   0.5696454251145529   0.8017179582594786   0.505608488956073   0.7693804886495247   0.8879550940134652   0.7938926295591058   0.4364971828254552   0.2153879916952374   0.7823943625603527   0.9105115172040619   0.7894930118246725   0.14361935358475061   0.8544570844032908   0.2798814999342015   0.3107920609739793   0.8392038808152767   0.8724695076685853   0.8880769507491584   0.07631679566260752   0.6461994557313486   0.3439481464371361   0.7054571914071167   0.25315429684789625   0.23750159300863902   0.7743027213225833   0.9037392331476382   0.7475458078918232   0.4681211043591143   0.8863476273091181   0.1098466035885324   0.31104862506636805   0.25273311266387694   0.1039532647487654   0.19933508638447056   0.5215556132416955   0.10911375907912632   0.24949618034547458   0.919453586450269   0.2107635522677162   0.26990987826384955   0.3770266726768893   0.03137663570111068   0.13444675660510869   0.6237104225325009   0.03307852623975316   0.32591944429399394   0.8812924597572124   0.3862088295238619   0.2587758049171699   0.4221802111463558   0.13374665186538923   0.9180877251647476
0.37242817760805186   0.31233360755782336   0.8226980267990212   0.6653546125008706   0.26847491285928643   0.11299852117335281   0.3011424135573257   0.5562408534217443   0.01897873251381186   0.1935449347230838   0.09037886128960945   0.2863309751578948   0.6419520598369226   0.1621682990219731   0.9559321046845007   0.6626205526253939   0.6088735335971694   0.8362488547279792   0.07463964492728833   0.27641172310153195   0.35009772867999955   0.4140686435816234   0.9408929930618991   0.3583239979367844   0.9776695510719478   0.10173503602380002   0.11819496626287791   0.6929693854359138   0.7091946382126613   0.9887365148504472   0.8170525527055522   0.13672853201416946   0.6902159056988494   0.7951915801273635   0.7266736914159428   0.8503975568562747   0.048263845861926793   0.6330232811053903   0.770741586731442   0.1877770042308808   0.43939031226475733   0.7967744263774111   0.6961019418041537   0.9113652811293488   0.0892925835847578   0.38270578279578776   0.7552089487422545   0.5530412831925644   0.11162303251281011   0.2809707467719877   0.6370139824793767   0.8600718977566507   0.4024283943001489   0.2922342319215405   0.8199614297738244   0.7233433657424813   0.7122124886012995   0.49704265179417706   0.09328773835788162   0.8729458088862065   0.6639486427393727   0.8640193706887868   0.32254615162643957   0.6851688046553258
0.22455833047461532   0.06724494431137565   0.6264442098222859   0.7738035235259769   0.13526574688985749   0.6845391615155879   0.8712352610800314   0.2207622403334125   0.02364271437704739   0.40356841474360017   0.23422127860065467   0.3606903425767618   0.6212143200768986   0.11133418282205969   0.41425984882683026   0.6373469768342805   0.9090018314755991   0.6142915310278826   0.32097211046894863   0.764401167948074   0.24505318873622642   0.7502721603390958   0.9984259588425091   0.07923236329274826   0.020494858261611102   0.6830272160277202   0.37198174902022313   0.3054288397667713   0.8852291113717536   0.9984880545121323   0.5007464879401918   0.08466659943335883   0.8615863969947062   0.5949196397685321   0.26652520933953716   0.7239762568565971   0.24037207691780768   0.4835854569464724   0.8522653605127068   0.08662928002231643   0.3313702454422086   0.8692939259185898   0.5312932500437583   0.3222281120742424   0.0863170567059822   0.11902176557949397   0.5328672912012492   0.24299574878149416   0.06582219844437111   0.4359945495517738   0.1608855421810261   0.9375669090147228   0.1805930870726175   0.4375064950396415   0.6601390542408343   0.852900309581364   0.31900669007791127   0.8425868552711094   0.39361384490129714   0.12892405272476698   0.07863461316010359   0.359001398324637   0.5413484843885902   0.042294772702450564
0.747264367717895   0.4897074724060472   0.010055234344831956   0.7200666606282081   0.6609473110119127   0.3706857068265532   0.4771879431435827   0.477070911846714   0.5951251125675416   0.9346911572747795   0.31630240096255663   0.5395040028319912   0.4145320254949242   0.49718466223513796   0.6561633467217224   0.6866036932506272   0.0955253354170129   0.6545978069640286   0.2625495018204252   0.5576796405258602   0.016890722256909303   0.2955964086393915   0.721201017431835   0.5153848678234096   0.26962635453901435   0.8058889362333443   0.711145783087003   0.7953182071952014   0.6086790435271016   0.4352032294067911   0.23395783994342031   0.31824729534848745   0.013553930959559866   0.5005120721320117   0.9176554389808637   0.7787432925164963   0.5990219054646357   0.0033274098968737544   0.26149209225914133   0.09213959926586911   0.5034965700476228   0.3487296029328452   0.9989425904387161   0.534459958740009   0.4866058477907135   0.05313319429345367   0.2777415730068811   0.019075090916599313   0.21697949325169916   0.24724425806010933   0.5665957899198781   0.22375688372139788   0.6083004497245976   0.8120410286533182   0.3326379499764578   0.9055095883729104   0.5947465187650377   0.3115289565213065   0.4149825109955941   0.12676629585641414   0.9957246133004021   0.3082015466244327   0.15349041873645275   0.03462669659054505
0.4922280432527793   0.9594719436915875   0.15454782829773664   0.5001667378505361   0.005622195462065797   0.9063387493981339   0.8768062552908555   0.4810916469339368   0.7886427022103666   0.6590944913380246   0.3102104653709774   0.25733476321253895   0.18034225248576902   0.8470534626847064   0.9775725153945196   0.35182517483962855   0.5855957337207313   0.5355245061633999   0.5625900043989256   0.2250588789832144   0.5898711204203292   0.22732295953896708   0.4090995856624728   0.19043218239266932   0.09764307716754994   0.2678510158473796   0.2545517573647362   0.6902654445421332   0.09202088170548414   0.3615122664492457   0.37774550207388063   0.2091737976081964   0.3033781794951175   0.7024177751112212   0.06753503670290321   0.9518390343956574   0.12303592700934847   0.8553643124265148   0.08996252130838357   0.6000138595560289   0.5374401932886173   0.319839806263115   0.5273725169094581   0.37495498057281457   0.947569072868288   0.09251684672414791   0.11827293124698524   0.18452279818014522   0.849925995700738   0.8246658308767684   0.8637211738822491   0.494257353638012   0.757905113995254   0.46315356442752265   0.4859756718083685   0.2850835560298156   0.4545269345001364   0.7607357893163015   0.41844063510546525   0.33324452163415813   0.3314910074907879   0.9053714768897866   0.3284781137970817   0.7332306620781293
0.7940508142021707   0.5855316706266717   0.8011055968876236   0.3582756815053147   0.8464817413338828   0.4930148239025237   0.6828326656406384   0.17375288332516947   0.9965557456331448   0.6683489930257553   0.8191114917583893   0.6794955296871574   0.2386506316378908   0.20519542859823273   0.33313581995002084   0.3944119736573419   0.7841236971377544   0.4444596392819312   0.9146951848445556   0.0611674520231837   0.45263268964696646   0.5390881623921446   0.586217071047474   0.3279367899450545   0.6585818754447957   0.953556491765473   0.7851114741598503   0.9696611084397397   0.812100134110913   0.46054166786294926   0.10227880851921191   0.7959082251145703   0.8155443884777682   0.7921926748371939   0.2831673167608226   0.11641269542741285   0.5768937568398774   0.5869972462389612   0.9500314968108017   0.722000721770071   0.7927700597021231   0.14253760695702994   0.035336311966246085   0.6608332697468873   0.34013737005515665   0.6034494445648854   0.44911924091877214   0.3328964798018328   0.6815554946103609   0.6498929527994124   0.6640077667589218   0.363235371362093   0.869455360499448   0.1893512849364631   0.5617289582397099   0.5673271462475227   0.05391097202167978   0.3971586100992692   0.27856164147888735   0.45091445082010984   0.47701721518180235   0.8101613638603081   0.3285301446680856   0.7289137290500388
0.6842471554796793   0.6676237569032781   0.2931938327018395   0.06808045930315158   0.34410978542452264   0.06417431233839281   0.8440745917830674   0.7351839795013188   0.6625542908141617   0.41428135953898043   0.1800668250241456   0.37194860813922576   0.7930989303147137   0.22493007460251732   0.6183378667844357   0.804621461891703   0.739187958293034   0.8277714645032481   0.33977622530554835   0.3537070110715932   0.26217074311123156   0.017610100642940003   0.011246080637462703   0.6247932820215544   0.5779235876315523   0.34998634373966186   0.7180522479356232   0.5567128227184027   0.2338138022070297   0.28581203140126904   0.8739776561525557   0.821528843217084   0.571259511392868   0.8715306718622886   0.6939108311284102   0.4495802350778582   0.7781605810781542   0.6466005972597713   0.07557296434397452   0.6449587731861552   0.03897262278512035   0.8188291327565232   0.7357967390384262   0.291251762114562   0.7768018796738888   0.8012190321135833   0.7245506584009634   0.6664584800930077   0.19887829204233645   0.45123268837392133   0.006498410465340325   0.10974565737460493   0.9650644898353068   0.1654206569726523   0.13252075431278457   0.28821681415752093   0.3938049784424388   0.2938899851103637   0.43860992318437436   0.8386365790796627   0.6156443973642846   0.6472893878505924   0.3630369588403999   0.1936778058935075
0.5766717745791642   0.8284602550940692   0.6272402198019736   0.9024260437789455   0.7998698949052754   0.02724122298048595   0.9026895614010102   0.23596756368593783   0.600991602862939   0.5760085346065646   0.8961911509356698   0.1262219063113329   0.6359271130276322   0.4105878776339123   0.7636703966228853   0.838005092153812   0.2421221345851934   0.11669789252354862   0.3250604734385109   0.9993685130741493   0.6264777372209089   0.46940850467295625   0.9620235145981111   0.8056907071806417   0.049805962641744715   0.6409482495788871   0.3347832947961374   0.9032646634016963   0.24993606773646931   0.6137070265984012   0.43209373339512724   0.6672970997157585   0.6489444648735303   0.037698491991836516   0.5359025824594574   0.5410751934044256   0.013017351845898145   0.6271106143579243   0.772232185836572   0.7030701012506135   0.7708952172607048   0.5104127218343756   0.4471717123980612   0.7037015881764643   0.14441748003979585   0.04100421716141937   0.48514819779995016   0.8980108809958225   0.09461151739805114   0.4000559675825323   0.15036490300381275   0.9947462175941263   0.8446754496615818   0.7863489409841312   0.7182711696086855   0.32744911787836783   0.1957309847880515   0.7486504489922947   0.18236858714922816   0.7863739244739423   0.18271363294215334   0.12153983463437046   0.41013640131265605   0.08330382322332874
0.4118184156814486   0.6111271127999949   0.9629646889145949   0.37960223504686447   0.26740093564165274   0.5701228956385755   0.4778164911146447   0.481591354051042   0.1727894182436016   0.17006692805604318   0.32745158811083197   0.4868451364569157   0.32811396858201974   0.38371798707191196   0.6091804185021464   0.15939601857854788   0.13238298379396826   0.6350675380796174   0.4268118313529183   0.3730220941046056   0.9496693508518149   0.5135277034452468   0.016675430040262233   0.28971827088127683   0.5378509351703663   0.902400590645252   0.053710741125667386   0.9101160358344124   0.27044999952871357   0.3322776950066765   0.5758942500110227   0.4285246817833704   0.09766058128511194   0.1622107669506333   0.24844266190019074   0.9416795453264547   0.7695466127030922   0.7784927798787213   0.6392622433980444   0.7822835267479068   0.6371636289091239   0.14342524179910401   0.21245041204512605   0.4092614326433012   0.687494278057309   0.6298975383538572   0.19577498200486382   0.11954316176202442   0.1496433428869427   0.7274969477086052   0.14206424087919645   0.20942712592761206   0.8791933433582292   0.3952192527019287   0.5661699908681738   0.7809024441442416   0.7815327620731172   0.2330084857512954   0.317727328967983   0.8392228988177869   0.011986149370025012   0.45451570587257406   0.6784650855699387   0.05693937206988009
0.3748225204609011   0.3110904640734701   0.46601467352481263   0.6476779394265788   0.6873282424035921   0.6811929257196129   0.2702396915199488   0.5281347776645544   0.5376848995166494   0.9536959780110077   0.12817545064075234   0.3187076517369424   0.6584915561584203   0.558476725309079   0.5620054597725785   0.5378052075927007   0.8769587940853031   0.3254682395577836   0.2442781308045956   0.6985823087749138   0.864972644715278   0.8709525336852095   0.5658130452346569   0.6416429367050337   0.49015012425437693   0.5598620696117395   0.09979837170984432   0.9939649972784549   0.8028218818507848   0.8786691438921266   0.8295586801898955   0.4658302196139005   0.26513698233413546   0.9249731658811189   0.7013832295491432   0.1471225678769581   0.6066454261757152   0.3664964405720399   0.1393777697765646   0.6093173602842574   0.7296866320904121   0.0410282010142563   0.895099638971969   0.9107350515093435   0.864713987375134   0.1700756673290468   0.32928659373731206   0.26909211480430983   0.3745638631207571   0.6102135977173073   0.22948822202746774   0.27512711752585495   0.5717419812699722   0.7315444538251809   0.39992954183757223   0.8092968979119545   0.3066049989358368   0.806571287944062   0.698546312288429   0.6621743300349964   0.6999595727601217   0.44007484737202207   0.5591685425118644   0.05285696975073903
0.9702729406697095   0.39904664635776577   0.6640689035398954   0.14212191824139545   0.10555895329457543   0.22897097902871896   0.3347823098025834   0.8730298034370856   0.7309950901738184   0.6187573813114116   0.10529408777511562   0.5979026859112306   0.15925310890384609   0.8872129274862308   0.7053645459375434   0.7886057879992762   0.8526481099680092   0.08064163954216887   0.006818233649114364   0.1264314579642797   0.15268853720788766   0.6405667921701468   0.4476496911372499   0.07357448821354068   0.18241559653817815   0.24152014581238104   0.7835807875973545   0.9314525699721452   0.07685664324360272   0.012549166783662085   0.4487984777947711   0.05842276653505962   0.3458615530697844   0.39379178547225047   0.34350439001965544   0.460520080623829   0.18660844416593833   0.5065788579860196   0.6381398440821121   0.6719142926245528   0.3339603341979291   0.4259372184438508   0.6313216104329977   0.5454828346602731   0.1812717969900414   0.785370426273704   0.18367191929574778   0.47190834644673246   0.9988562004518633   0.543850280461323   0.40009113169839333   0.5404557764745872   0.9219995572082605   0.5313011136776609   0.9512926539036223   0.48203300993952763   0.5761380041384762   0.13750932820541037   0.6077882638839668   0.021512929315698637   0.3895295599725378   0.6309304702193907   0.9696484198018547   0.34959863669114577
0.055569225774608724   0.2049932517755399   0.338326809368857   0.8041158020308726   0.8742974287845673   0.41962282550183594   0.15465489007310923   0.3322074555841401   0.8754412283327041   0.8757725450405129   0.7545637583747159   0.7917516791095529   0.9534416711244436   0.34447143136285213   0.8032711044710937   0.3097186691700253   0.37730366698596746   0.20696210315744173   0.19548284058712692   0.2882057398543266   0.9877741070134296   0.576031632938051   0.22583442078527222   0.9386071031631809   0.932204881238821   0.3710383811625111   0.8875076114164152   0.13449130113230826   0.057907452454253605   0.9514155556606751   0.7328527213433059   0.8022838455481681   0.18246622412154953   0.07564301062016221   0.97828896296859   0.01053216643861524   0.22902455299710597   0.7311715792573101   0.17501785849749632   0.70081349726859   0.8517208860111385   0.5242094760998683   0.9795350179103693   0.41260775741426337   0.8639467789977089   0.9481778431618173   0.7537005971250972   0.4740006542510825   0.9317418977588879   0.5771394619993062   0.866192985708682   0.3395093531187743   0.8738344453046344   0.6257239063386311   0.133340264365376   0.5372255075706062   0.6913682211830848   0.5500808957184689   0.15505130139678597   0.526693341131991   0.46234366818597883   0.8189093164611587   0.9800334428992896   0.825879843863401
0.6106227821748403   0.2946998403612904   0.0004984249889202434   0.41327208644913754   0.7466760031771315   0.346521997199473   0.24679782786382307   0.939271432198055   0.8149341054182434   0.7693825352001668   0.3806048421551411   0.5997620790792807   0.9410996601136091   0.14365862886153571   0.2472645777897651   0.06253657150867456   0.2497314389305243   0.5935777331430669   0.09221327639297913   0.5358432303766836   0.7873877707445455   0.7746684166819081   0.11217983349368948   0.7099633865132827   0.17676498856970516   0.4799685763206178   0.11168140850476925   0.2966913000641451   0.43008898539257373   0.1334465791211448   0.8648835806409462   0.3574198678660901   0.6151548799743303   0.364064043920978   0.48427873848580505   0.7576577887868093   0.6740552198607211   0.22040541505944228   0.23701416069603998   0.6951212172781348   0.4243237809301969   0.6268276819163754   0.14480088430306085   0.1592779869014512   0.6369360101856515   0.8521592652344673   0.03262105080937135   0.4493146003881685   0.4601710216159463   0.37219068891384943   0.9209396423046021   0.1526233003240234   0.03008203622337253   0.23874410979270463   0.05605606166365593   0.7952034324579332   0.41492715624904225   0.8746800658717266   0.5717773231778509   0.03754564367112391   0.740871936388321   0.6542746508122843   0.33476316248181087   0.3424244263929891
0.31654815545812415   0.027446968895908936   0.18996227817875005   0.1831464394915379   0.6796121452724727   0.17528770366144172   0.1573412273693787   0.7338318391033694   0.21944112365652643   0.8030970147475923   0.23640158506477657   0.581208538779346   0.18935908743315388   0.5643529049548877   0.18034552340112064   0.7860051063214126   0.7744319311841117   0.689672839083161   0.6085682002232697   0.7484594626502887   0.03355999479579062   0.03539818827087672   0.27380503774145887   0.4060350362572997   0.7170118393376664   0.007951219374967783   0.08384275956270884   0.2228885967657618   0.03739969406519377   0.832663515713526   0.9265015321933302   0.4890567576623924   0.8179585704086674   0.029566500965933783   0.6900999471285536   0.9078482188830465   0.6285994829755135   0.4652135960110461   0.509754423727433   0.12184311256163383   0.8541675517914018   0.775540756927885   0.9011862235041631   0.37338364991134504   0.8206075569956112   0.7401425686570083   0.6273811857627043   0.9673486136540453   0.1035957176579447   0.7321913492820405   0.5435384261999954   0.7444600168882836   0.06619602359275094   0.8995278335685145   0.6170368940066653   0.25540325922589113   0.24823745318408358   0.8699613326025807   0.9269369468781117   0.3475550403428446   0.6196379702085701   0.40474773659153457   0.4171825231506787   0.2257119277812108
0.7654704184171683   0.6292069796636495   0.5159962996465156   0.8523282778698658   0.9448628614215572   0.8890644110066411   0.8886151138838113   0.8849796642158203   0.8412671437636124   0.15687306172460058   0.3450766876838159   0.14051964732753677   0.7750711201708615   0.25734522815608607   0.7280397936771507   0.8851163881016456   0.5268336669867779   0.3873838955535054   0.801102846799039   0.537561347758801   0.9071956967782078   0.9826361589619708   0.3839203236483602   0.3118494199775902   0.14172527836103946   0.35342917929832124   0.8679240240018447   0.4595211421077245   0.19686241693948234   0.4643647682916801   0.9793089101180333   0.5745414778919041   0.35559527317586986   0.3074917065670795   0.6342322224342174   0.4340218305643674   0.5805241530050084   0.05014647841099342   0.9061924287570667   0.5489054424627218   0.05369048601823047   0.662762582857488   0.10508958195802784   0.011344094703920712   0.14649478924002268   0.6801264238955173   0.7211692583096676   0.6994946747263305   0.0047695108789832085   0.326697244597196   0.8532452343078231   0.23997353261860602   0.8079070939395009   0.8623324763055159   0.8739363241897897   0.6654320547267019   0.45231182076363097   0.5548407697384364   0.23970410175557233   0.2314102241623345   0.8717876677586226   0.504694291327443   0.33351167299850554   0.6825047816996128
0.8180971817403921   0.8419317084699549   0.2284220910404777   0.6711606869956921   0.6716023925003695   0.16180528457443766   0.50725283273081   0.9716660122693616   0.6668328816213862   0.8351080399772416   0.6540075984229871   0.7316924796507556   0.8589257876818853   0.9727755636717257   0.7800712742331973   0.06626042492405368   0.40661396691825435   0.4179347939332893   0.540367172477625   0.8348502007617191   0.5348262991596318   0.9132405026058463   0.20685549947911944   0.15234541906210639   0.7167291174192396   0.07130879413589142   0.9784334084386418   0.4811847320664143   0.045126724918870174   0.9095035095614538   0.4711805757078317   0.5095187197970528   0.37829384329748394   0.07439546958421213   0.8171729772848446   0.7778262401462972   0.5193680556155986   0.1016199059124864   0.037101703051647346   0.7115658152222435   0.1127540886973442   0.6836851119791971   0.49673453057402234   0.8767156144605243   0.5779277895377124   0.7704446093733508   0.28987903109490293   0.724370195398418   0.8611986721184728   0.6991358152374594   0.3114456226562612   0.24318546333200364   0.8160719471996026   0.7896323056760056   0.8402650469484295   0.7336667435349509   0.4377781039021187   0.7152368360917934   0.02309206966358483   0.9558405033886538   0.9184100482865202   0.6136169301793071   0.9859903666119375   0.2442746881664103
0.8056559595891759   0.92993181820011   0.4892558360379151   0.367559073705886   0.2277281700514635   0.1594872088267592   0.19937680494301221   0.6431888783074681   0.36652949793299067   0.4603513935892999   0.887931182286751   0.4000034149754644   0.5504575507333881   0.6707190879132943   0.047666135338321564   0.6663366714405135   0.11267944683126938   0.9554822518215008   0.02457406567473673   0.7104961680518597   0.19426939854474926   0.3418653216421938   0.038583699062799244   0.46622147988544943   0.3886134389555733   0.41193350344208385   0.5493278630248841   0.09866240617956346   0.16088526890410984   0.25244629461532464   0.34995105808187194   0.45547352787209544   0.7943557709711191   0.7920949010260248   0.4620198757951209   0.055470112896631035   0.24389822023773106   0.12137581311273045   0.4143537404567993   0.38913344145611756   0.13121877340646168   0.16589356129122962   0.3897796747820626   0.6786372734042578   0.9369493748617125   0.8240282396490358   0.3511959757192633   0.21241579351880846   0.5483359359061392   0.412094736206952   0.8018681126943792   0.113753387339245   0.3874506670020293   0.15964844159162736   0.4519170546125073   0.6582798594671496   0.5930948960309101   0.36755354056560263   0.9898971788173865   0.6028097465705186   0.3491966757931791   0.24617772745287217   0.5755434383605871   0.21367630511440097
0.21797790238671738   0.08028416616164256   0.18576376357852456   0.5350390317101431   0.28102852752500496   0.25625592651260676   0.8345677878592612   0.32262323819133465   0.7326925916188658   0.8441611903056547   0.03269967516488201   0.20886985085208962   0.34524192461683656   0.6845127487140273   0.5807826205523747   0.55058999138494   0.7521470285859264   0.31695920814842476   0.5908854417349882   0.9477802448144215   0.4029503527927473   0.07078148069555258   0.015342003374401147   0.7341039397000205   0.18497245040602991   0.99049731453391   0.8295782397958766   0.19906490798987744   0.903943922881025   0.7342413880213032   0.9950104519366154   0.8764416697985428   0.17125133126215913   0.8900801977156485   0.9623107767717334   0.6675718189464531   0.8260094066453226   0.20556744900162113   0.38152815621935865   0.11698182756151312   0.07386237805939619   0.8886082408531963   0.7906427144843704   0.16920158274709163   0.6709120252666488   0.8178267601576438   0.7753007111099692   0.4350976430470711   0.48593957486061895   0.8273294456237338   0.9457224713140927   0.23603273505719366   0.581995651979594   0.09308805760243048   0.9507120193774773   0.35959106525865087   0.4107443207174349   0.20300785988678197   0.9884012426057439   0.6920192463121977   0.5847349140721123   0.9974404108851608   0.6068730863863853   0.5750374187506846
0.5108725360127161   0.10883217003196446   0.8162303719020149   0.40583583600359296   0.8399605107460673   0.29100540987432066   0.04092966079204557   0.9707381929565219   0.35402093588544825   0.46367596425058694   0.09520718947795291   0.7347054578993282   0.7720252839058543   0.37058790664815644   0.14449517010047563   0.3751143926406773   0.3612809631884194   0.16758004676137447   0.15609392749473175   0.6830951463284796   0.7765460491163071   0.17013963587621364   0.5492208411083466   0.10805772757779503   0.26567351310359105   0.06130746584424917   0.7329904692063317   0.702221891574202   0.4257130023575238   0.7703020559699285   0.6920608084142862   0.7314836986176801   0.07169206647207553   0.3066260917193416   0.5968536189363333   0.996778240718352   0.29966678256622126   0.9360381850711852   0.4523584488358576   0.6216638480776747   0.9383858193778019   0.7684581383098107   0.29626452134112585   0.938568701749195   0.16183977026149468   0.5983185024335971   0.7470436802327793   0.8305109741714001   0.8961662571579037   0.5370110365893479   0.014053211026447604   0.12828908259719798   0.4704532548003798   0.7667089806194194   0.32199240261216144   0.3968053839795178   0.39876118832830426   0.4600828889000778   0.7251387836758282   0.4000271432611658   0.09909440576208303   0.5240447038288927   0.2727803348399706   0.7783632951834911
0.1607085863842812   0.755586565519082   0.9765158134988448   0.8397945934342961   0.9988688161227866   0.1572680630854849   0.22947213326606547   0.009283619262895967   0.10270255896488291   0.620257026496137   0.21541892223961787   0.8809945366656979   0.6322493041645031   0.8535480458767176   0.8934265196274565   0.4841891526861802   0.2334881158361988   0.3934651569766398   0.1682877359516282   0.08416200942501438   0.13439371007411577   0.8694204531477471   0.8955074011116575   0.3057987142415233   0.9736851236898345   0.11383388762866513   0.9189915876128127   0.46600412080722725   0.9748163075670481   0.9565658245431802   0.6895194543467473   0.4567205015443313   0.8721137486021652   0.3363087980470432   0.47410053210712944   0.5757259648786333   0.23986444443766203   0.4827607521703256   0.580674012479673   0.09153681219245313   0.006376328601463221   0.08929559519368582   0.4123862765280449   0.00737480276743876   0.8719826185273475   0.21987514204593872   0.5168788754163873   0.7015760885259155   0.8982974948375129   0.10604125441727358   0.5978872878035746   0.23557196771868824   0.9234811872704649   0.14947542987409337   0.9083678334568273   0.778851466174357   0.05136743866829974   0.8131666318270502   0.4342673013496978   0.20312550129572365   0.8115029942306378   0.3304058796567246   0.8535932888700247   0.11158868910327051
0.8051266656291745   0.24111028446303873   0.4412070123419799   0.10421388633583174   0.9331440471018271   0.021235142417100027   0.9243281369255926   0.40263779780991626   0.034846552264314164   0.9151938879998265   0.32644084912201804   0.16706583009122802   0.1113653649938493   0.765718458125733   0.4180730156651908   0.3882143639168711   0.05999792632554956   0.952551826298683   0.983805714315493   0.18508886262114743   0.24849493209491186   0.6221459466419583   0.13021242544546827   0.07350017351787692   0.44336826646573735   0.38103566217891965   0.6890054131034884   0.9692862871820451   0.5102242193639103   0.3598005197618196   0.7646772761778958   0.566648489372129   0.47537766709959617   0.44460663176199317   0.43823642705587773   0.3995826592809009   0.36401230210574687   0.6788881736362601   0.020163411390686926   0.011368295364029824   0.3040143757801973   0.7263363473375771   0.036357697075193915   0.8262794327428824   0.05551944368528544   0.10419040069561879   0.9061452716297257   0.7527792592250054   0.612151177219548   0.7231547385166992   0.2171398585262373   0.7834929720429603   0.10192695785563778   0.36335421875487955   0.4524625823483415   0.2168444826708314   0.6265492907560416   0.9187475869928864   0.014226155292463794   0.8172618233899305   0.2625369886502948   0.23985941335662633   0.9940627439017768   0.8058935280259006
0.9585226128700975   0.5135230660190492   0.957705046826583   0.9796140952830182   0.903003169184812   0.4093326653234304   0.05155977519685729   0.2268348360580128   0.29085199196526396   0.6861779268067312   0.83441991667062   0.4433418640150525   0.1889250341096262   0.3228237080518516   0.38195733432227846   0.2264973813442211   0.5623757433535845   0.40407612105896523   0.36773117902981467   0.4092355579542906   0.29983875470328974   0.16421670770233893   0.3736684351280378   0.6033420299283899   0.34131614183319225   0.6506936416832897   0.41596338830145485   0.6237279346453717   0.4383129726483802   0.24136097635985937   0.36440361310459757   0.3968930985873589   0.14746098068311622   0.5551830495531281   0.5299836964339776   0.9535512345723064   0.9585359465734901   0.23235934150127652   0.14802636211169912   0.7270538532280852   0.39616020321990547   0.8282832204423113   0.7802951830818844   0.3178182952737947   0.09632144851661573   0.6640665127399724   0.4066267479538466   0.7144762653454048   0.7550053066834235   0.01337287105668262   0.9906633596523918   0.09074833070003305   0.31669233403504327   0.7720118946968233   0.6262597465477943   0.6938552321126742   0.16923135335192704   0.21682884514369508   0.09627605011381665   0.7403039975403678   0.210695406778437   0.9844695036424186   0.9482496880021175   0.013250144312282473
0.8145352035585315   0.1561862832001073   0.1679545049202331   0.6954318490384878   0.7182137550419158   0.49211977046013494   0.7613277569663864   0.9809555836930831   0.9632084483584923   0.47874689940345233   0.7706643973139947   0.89020725299305   0.646516114323449   0.7067350047066291   0.14440465076620046   0.19635202088037587   0.477284760971522   0.489906159562934   0.0481286006523838   0.4560480233400081   0.266589354193085   0.5054366559205153   0.09987891265026626   0.44279787902772566   0.4520541506345535   0.3492503727204081   0.9319244077300332   0.7473660299892378   0.7338403955926377   0.8571306022602732   0.1705966507636467   0.7664104462961547   0.7706319472341454   0.3783837028568209   0.399932253449652   0.8762031933031047   0.1241158329106963   0.6716486981501918   0.25552760268345154   0.6798511724227289   0.6468310719391743   0.18174253858725783   0.20739900203106776   0.22380314908272073   0.3802417177460893   0.6763058826667424   0.10752008938080151   0.7810052700549951   0.9281875671115358   0.32705550994633437   0.17559568165076836   0.033639240065757234   0.1943471715188981   0.46992490768606116   0.004999030887121662   0.26722879376960246   0.4237152242847528   0.0915412048292403   0.6050667774374696   0.39102560046649776   0.29959939137405645   0.4198925066790485   0.3495391747540181   0.7111744280437688
0.6527683194348821   0.23814996809179065   0.14214017272295032   0.48737127896104815   0.2725266016887929   0.5618440854250482   0.034620083342148805   0.7063660089060531   0.34433903457725706   0.23478857547871385   0.8590244016913805   0.6727267688402958   0.14999186305835896   0.7648636677926527   0.8540253708042588   0.4054979750706934   0.7262766387736062   0.6733224629634124   0.24895859336678913   0.014472374604195641   0.42667724739954976   0.2534299562843639   0.8994194186127711   0.30329794656042675   0.7739089279646676   0.015279988192573217   0.7572792458898208   0.8159266675993786   0.5013823262758748   0.45343590276752505   0.7226591625476719   0.10956065869332551   0.15704329169861764   0.21864732728881117   0.8636347608562915   0.4368338898530297   0.00705142864025868   0.4537836594961585   0.009609390052032712   0.031335914782336285   0.2807747898666525   0.7804611965327461   0.7606507966852436   0.016863540178140644   0.8540975424671027   0.5270312402483823   0.8612313780724725   0.7135655936177139   0.08018861450243515   0.5117512520558091   0.10395213218265177   0.8976389260183353   0.5788062882265604   0.058315349288284045   0.38129296963497983   0.7880782673250097   0.4217629965279428   0.8396680219994729   0.5176582087786883   0.3512443774719801   0.41471156788768415   0.38588436250331437   0.5080488187266556   0.31990846268964385
0.13393677802103165   0.6054231659705682   0.747398022041412   0.30304492251150317   0.2798392355539289   0.07839192572218592   0.8861666439689395   0.5894793288937893   0.19965062105149375   0.5666406736663768   0.7822145117862878   0.691840402875454   0.6208443328249333   0.5083253243780929   0.40092154215130793   0.9037621355504442   0.1990813362969905   0.66865730237862   0.8832633333726196   0.552517758078464   0.7843697684093064   0.2827729398753056   0.375214514645964   0.23260929538882025   0.6504329903882747   0.6773497739047374   0.627816492604552   0.9295643728773171   0.3705937548343458   0.5989578481825515   0.7416498486356125   0.3400850439835278   0.17094313378285209   0.032317174516174614   0.9594353368493247   0.6482446411080738   0.5500988009579187   0.5239918501380818   0.5585137946980168   0.7444825055576295   0.35101746466092826   0.8553345477594618   0.6752504613253971   0.19196474747916548   0.5666476962516218   0.5725616078841562   0.3000359466794331   0.9593554520903452   0.9162147058633471   0.8952118339794188   0.6722194540748812   0.029791079213028173   0.5456209510290012   0.2962539857968674   0.9305696054392687   0.6897060352295004   0.3746778172461492   0.2639368112806928   0.971134268589944   0.04146139412142664   0.8245790162882304   0.739944961142611   0.4126204738919273   0.29697888856379706
0.4735615516273022   0.8846104133831492   0.7373700125665302   0.10501414108463158   0.9069138553756804   0.31204880549899283   0.43733406588709706   0.14565868899428636   0.9906991495123333   0.416836971519574   0.765114611812216   0.11586760978125818   0.445078198483332   0.12058298572270655   0.8345450063729472   0.4261615745517578   0.07040038123718284   0.8566461744420137   0.8634107377830031   0.3847001804303311   0.24582136494895243   0.11670121329940275   0.45079026389107585   0.08772129186653406   0.7722598133216503   0.23209079991625362   0.7134202513245457   0.9827071507819025   0.8653459579459699   0.9200419944172608   0.2760861854374486   0.8370484617876162   0.8746468084336366   0.5032050228976868   0.5109715736252327   0.721180852006358   0.4295686099503046   0.3826220371749802   0.6764265672522856   0.29501927745460016   0.35916822871312176   0.5259758627329665   0.8130158294692823   0.910319097024269   0.11334686376416936   0.40927464943356373   0.3622255655782065   0.822597805157735   0.3410870504425191   0.17718384951731012   0.6488053142536608   0.8398906543758325   0.4757410924965492   0.25714185510004933   0.3727191288162122   0.0028421925882163783   0.6010942840629125   0.7539368322023625   0.8617475551909796   0.28166134058185843   0.17152567411260794   0.3713147950273823   0.185320987938694   0.9866420631272582
0.8123574453994862   0.8453389322944158   0.37230515846941165   0.07632296610298922   0.6990105816353168   0.4360642828608521   0.010079592891205162   0.25372516094525427   0.3579235311927977   0.258880433343542   0.36127427863754435   0.4138345065694217   0.8821824386962485   0.0017385782434926392   0.9885551498213321   0.4109923139812054   0.2810881546333359   0.2478017460411301   0.1268075946303526   0.12933097339934693   0.10956248052072798   0.8764869510137477   0.9414866066916586   0.14268891027208866   0.2972050351212418   0.031148018719331923   0.5691814482222469   0.06636594416909945   0.598194453485925   0.5950837358584798   0.5591018553310417   0.8126407832238453   0.24027092229312733   0.33620330251493785   0.19782757669349743   0.3988062766544235   0.35808848359687884   0.3344647242714452   0.20927242687216532   0.9878139626732181   0.07700032896354289   0.08666297823031512   0.08246483224181271   0.8584829892738711   0.9674378484428149   0.21017602721656736   0.1409782255501541   0.7157940790017825   0.6702328133215731   0.17902800849723544   0.5717967773279071   0.649428134832683   0.07203835983564807   0.5839442726387556   0.01269492199686539   0.8367873516088379   0.8317674375425208   0.24774097012381777   0.8148673453033679   0.4379810749544144   0.47367895394564197   0.9132762458523725   0.6055949184312026   0.45016711228119627
0.39667862498209905   0.8266132676220574   0.5231300861893899   0.5916841230073251   0.42924077653928416   0.6164372404054901   0.3821518606392358   0.8758900440055427   0.759007963217711   0.43740923190825465   0.8103550833113287   0.22646190917285963   0.6869696033820629   0.8534649592694991   0.7976601613144633   0.3896745575640218   0.8552021658395422   0.6057239891456813   0.9827928160110954   0.9516934826096074   0.38152321189390026   0.6924477432933087   0.3771978975798927   0.5015263703284111   0.9848445869118012   0.8658344756712513   0.8540678113905028   0.909842247321086   0.555603810372517   0.24939723526576113   0.47191595075126697   0.033952203315543314   0.796595847154806   0.8119880033575064   0.6615608674399382   0.8074902941426837   0.10962624377274305   0.9585230440880074   0.8639007061254751   0.4178157365786619   0.2544240779332009   0.3527990549423261   0.8811078901143797   0.4661222539690545   0.8729008660393006   0.6603513116490174   0.5039099925344871   0.9645958836406433   0.8880562791274994   0.7945168359777661   0.6498421811439843   0.054753636319557375   0.33245246875498236   0.545119600712005   0.17792623039271738   0.020801433004014058   0.5358566216001763   0.7331315973544985   0.516365362952779   0.21331113886133038   0.4262303778274333   0.7746085532664911   0.652464656827304   0.7954954022826685
0.1718062998942324   0.42180949832416503   0.7713567667129243   0.32937314831361403   0.2989054338549318   0.7614581866751476   0.2674467741784372   0.36477726467297067   0.4108491547274324   0.9669413506973815   0.6176045930344529   0.3100236283534133   0.07839668597245007   0.42182174998537647   0.43967836264173554   0.28922219534939925   0.5425400643722738   0.688690152630878   0.9233129996889565   0.07591105648806887   0.11630968654484049   0.9140815993643868   0.27084834286165244   0.2804156542054004   0.9445033866506081   0.4922721010402218   0.4994915761487282   0.9510425058917864   0.6455979527956762   0.7308139143650741   0.23204480197029095   0.5862652412188157   0.23474879806824386   0.7638725636676927   0.6144402089358381   0.2762416128654024   0.15635211209579378   0.3420508136823162   0.1747618462941025   0.9870194175160031   0.61381204772352   0.6533606610514383   0.251448846605146   0.9111083610279342   0.4975023611786795   0.7392790616870515   0.9806005037434935   0.6306927068225339   0.5529989745280715   0.24700696064682964   0.48110892759476537   0.6796502009307476   0.9074010217323952   0.5161930462817554   0.24906412562447444   0.09338495971193186   0.6726522236641513   0.7523204826140628   0.6346239166886364   0.8171433468465295   0.5163001115683575   0.41026966893174655   0.4598620703945339   0.8301239293305264
0.9024880638448376   0.7569090078803082   0.20841322378938792   0.9190155683025921   0.404985702666158   0.01762994619325684   0.22781272004589437   0.28832286148005815   0.8519867281380865   0.7706229855464272   0.7467037924511291   0.6086726605493106   0.9445857064056913   0.2544299392646717   0.49763966682665456   0.5152877008373787   0.27193348274154   0.502109456650609   0.8630157501380181   0.6981443539908493   0.7556333711731824   0.09183978771886242   0.4031536797434842   0.8680204246603229   0.8531453073283448   0.3349307798385541   0.1947404559540963   0.9490048563577309   0.44815960466218685   0.3173008336452973   0.9669277359082019   0.6606819948776727   0.5961728765241002   0.5466778480988701   0.2202239434570729   0.05200933432836207   0.6515871701184089   0.2922479088341984   0.7225842766304184   0.5367216334909833   0.379653687376869   0.7901384521835894   0.8595685264924002   0.838577279500134   0.6240203162036866   0.698298664464727   0.45641484674891597   0.9705568548398111   0.7708750088753418   0.3633678846261728   0.2616743907948197   0.02155199848208021   0.3227154042131549   0.04606705098087554   0.2947466548866177   0.3608700036044075   0.7265425276890546   0.49938920288200545   0.07452271142954482   0.30886066927604544   0.07495535757064568   0.2071412940478071   0.35193843479912645   0.7721390357850622
0.6953016701937768   0.4170028418642177   0.4923699083067263   0.9335617562849281   0.07128135399009014   0.7187041773994908   0.03595506155781031   0.9630049014451171   0.3004063451147484   0.3553362927733179   0.7742806707629907   0.9414529029630369   0.9776909409015935   0.30926924179244236   0.4795340158763729   0.5805828993586293   0.25114841321253883   0.8098800389104369   0.4050113044468281   0.2717222300825839   0.17619305564189316   0.6027387448626298   0.05307286964770161   0.49958319429752174   0.48089138544811644   0.1857359029984121   0.5607029613409753   0.5660214380125936   0.4096100314580263   0.4670317255989214   0.524747899783165   0.6030165365674766   0.10920368634327791   0.11169543282560351   0.7504672290201744   0.6615636336044398   0.13151274544168443   0.8024261910331612   0.2709332131438015   0.08098073424581047   0.8803643322291456   0.9925461521227242   0.8659219086969734   0.8092585041632265   0.7041712765872524   0.38980740726009444   0.8128490390492717   0.30967530986570485   0.223279891139136   0.20407150426168236   0.25214607770829645   0.7436538718531112   0.8136698596811097   0.7370397786627609   0.7273981779251314   0.1406373352856346   0.7044661733378318   0.6253443458371575   0.976930948904957   0.47907370168119484   0.5729534278961473   0.8229181548039962   0.7059977357611555   0.39809296743538436
0.6925890956670018   0.830372002681272   0.8400758270641822   0.5888344632721577   0.9884178190797493   0.44056459542117754   0.027226788014910366   0.2791591534064529   0.7651379279406133   0.23649309115949518   0.7750807103066139   0.5355052815533418   0.9514680682595037   0.49945331249673425   0.04768253238148248   0.3948679462677071   0.2470018949216719   0.8741089666595768   0.07075158347652542   0.9157942445865123   0.6740484670255246   0.05119081185558053   0.36475384771536984   0.5177012771511279   0.9814593713585228   0.22081880917430854   0.5246780206511877   0.9288668138789702   0.9930415522787736   0.780254213753131   0.49745123263627733   0.6497076604725173   0.2279036243381602   0.5437611225936358   0.7223705223296635   0.11420237891917553   0.2764355560786565   0.04430781009690163   0.6746879899481809   0.7193344326514685   0.029433661156984616   0.17019884343732483   0.6039364064716555   0.8035401880649561   0.35538519413146   0.1190080315817443   0.23918255875628566   0.2858389109138281   0.3739258227729372   0.8981892224074357   0.714504538105098   0.356972097034858   0.3808842704941637   0.11793500865430473   0.21705330546882062   0.7072644365623407   0.15298064615600349   0.5741738860606689   0.4946827831391572   0.5930620576431652   0.8765450900773469   0.5298660759637672   0.8199947931909762   0.8737276249916968
0.8471114289203624   0.3596672325264424   0.2160583867193207   0.07018743692674066   0.4917262347889023   0.24065920094469812   0.9768758279630351   0.7843485260129125   0.11780041201596513   0.34246997853726235   0.26237128985793706   0.42737642897805456   0.7369161415218014   0.22453496988295765   0.04531798438911646   0.7201119924157139   0.5839354953657979   0.6503610838222887   0.5506352012499592   0.12704993477254867   0.707390405288451   0.12049500785852152   0.730640408058983   0.2533223097808519   0.8602789763680887   0.7608277753320791   0.5145820213396624   0.18313487285411123   0.3685527415791863   0.520168574387381   0.5377061933766273   0.3987863468411987   0.25075232956322124   0.17769859585011863   0.2753349035186902   0.9714099178631441   0.5138361880414197   0.953163625967161   0.23001691912957373   0.25129792544743035   0.9299006926756218   0.30280254214487223   0.6793817178796144   0.12424799067488168   0.2225102873871708   0.18230753428635071   0.9487413098206314   0.8709256808940298   0.3622313110190822   0.4214797589542716   0.43415928848096913   0.6877908080399185   0.9936785694398959   0.9013111845668906   0.8964530951043418   0.28900446119871986   0.7429262398766746   0.7236125887167719   0.6211181915856516   0.3175945433355757   0.22909005183525483   0.7704489627496109   0.3911012724560779   0.06629661788814536
0.299189359159633   0.46764642060473877   0.7117195545764634   0.9420486272132637   0.07667907177246222   0.28533888631838805   0.762978244755832   0.07112294631923391   0.71444776075338   0.8638591273641164   0.3288189562748629   0.38333213827931534   0.7207691913134843   0.9625479427972259   0.43236586117052106   0.09432767708059547   0.9778429514368097   0.23893535408045388   0.8112476695848694   0.7767331337450197   0.7487528996015548   0.4684863913308429   0.4201463971287915   0.7104365158568744   0.44956354044192176   0.0008399707261041557   0.708426842552328   0.7683878886436107   0.37288446866945957   0.7155010844077161   0.945448597796496   0.6972649423243769   0.6584367079160794   0.8516419570435997   0.6166296415216331   0.31393280404506146   0.9376675166025953   0.8890940142463738   0.18426378035111213   0.219605126964466   0.9598245651657856   0.6501586601659199   0.3730161107662427   0.4428719932194462   0.2110716655642308   0.181672268835077   0.9528697136374512   0.7324354773625718   0.761508125122309   0.18083229810897283   0.24444287108512316   0.9640475887189611   0.38862365645284946   0.46533121370125674   0.2989942732886271   0.26678264639458427   0.73018694853677   0.6136892566576571   0.6823646317669939   0.9528498423495227   0.7925194319341747   0.7245952424112833   0.4981008514158818   0.7332447153850568
0.8326948667683891   0.07443658224536338   0.1250847406496391   0.29037272216561055   0.6216232012041584   0.8927643134102864   0.17221502701218788   0.5579372448030387   0.8601150760818493   0.7119320153013136   0.9277721559270647   0.5938896560840777   0.4714914196289998   0.2466008016000568   0.6287778826384376   0.3271070096894934   0.7413044710922299   0.6329115449423997   0.9464132508714437   0.3742571673399706   0.9487850391580551   0.9083163025311164   0.4483123994555619   0.6410124519549139   0.116090172389666   0.8338797202857531   0.3232276588059228   0.35063972978930324   0.49446697118550764   0.9411154068754667   0.15101263179373492   0.7927024849862645   0.6343518951036583   0.22918339157415313   0.22324047586667017   0.1988128289021868   0.1628604754746585   0.9825825899740963   0.5944625932282326   0.8717058192126934   0.42155600438242863   0.3496710450316966   0.6480493423567888   0.49744865187272275   0.4727709652243735   0.4413547425005802   0.19973694290122693   0.856436199917809   0.3566807928347075   0.6074750222148272   0.8765092840953042   0.5057964701285057   0.8622138216491999   0.6663596153393605   0.7254966523015692   0.7130939851422412   0.22786192654554152   0.43717622376520743   0.5022561764348991   0.5142811562400544   0.06500145107088301   0.4545936337911111   0.9077935832066665   0.6425753370273611
0.6434454466884544   0.10492258875941449   0.2597442408498777   0.14512668515463834   0.17067448146408087   0.6635678462588342   0.060007297948650756   0.2886904852368294   0.8139936886293734   0.056092824044007075   0.1834980138533466   0.7828940151083237   0.9517798669801735   0.3897332087046465   0.4580013615517774   0.06980002996608241   0.723917940434632   0.9525569849394391   0.9557451851168783   0.5555188737260279   0.658916489363749   0.497963351148328   0.047951601910211784   0.9129435366986669   0.015471042675294611   0.3930407623889135   0.7882073610603341   0.7678168515440286   0.8447965612112137   0.7294729161300793   0.7282000631116833   0.4791263663071992   0.030802872581840387   0.6733800920860722   0.5447020492583368   0.6962323511988755   0.07902300560166688   0.28364688338142563   0.08670068770655935   0.6264323212327931   0.3551050651670349   0.33108989844198655   0.13095550258968106   0.07091344750676516   0.6961885758032859   0.8331265472936585   0.08300390067946926   0.1579699108080983   0.6807175331279913   0.44008578490474504   0.29479653961913516   0.3901530592640698   0.8359209719167775   0.7106128687746658   0.5665964765074518   0.9110266929568707   0.8051180993349372   0.037232776688593594   0.021894427249115115   0.2147943417579951   0.7260950937332703   0.753585893307168   0.9351937395425558   0.588362020525202
0.37099002856623536   0.4224959948651814   0.8042382369528748   0.5174485730184368   0.6748014527629494   0.5893694475715229   0.7212343362734055   0.35947866221033853   0.9940839196349582   0.1492836626667778   0.4264377966542703   0.9693256029462688   0.15816294771818065   0.43867079389211205   0.8598413201468185   0.05829890998939815   0.3530448483832435   0.40143801720351846   0.8379468928977033   0.8435045682314031   0.6269497546499733   0.6478521238963505   0.9027531533551476   0.25514254770620104   0.25595972608373785   0.2253561290311691   0.09851491640227285   0.7376939746877642   0.5811582733207883   0.6359866814596462   0.3772805801288674   0.3782153124774256   0.5870743536858302   0.4867030187928684   0.950842783474597   0.40888970953115683   0.4289114059676495   0.04803222490075639   0.09100146332777866   0.3505907995417587   0.07586655758440598   0.646594207697238   0.25305457043007534   0.5070862313103557   0.44891680293443276   0.9987420838008875   0.35030141707492773   0.25194368360415464   0.19295707685069494   0.7733859547697183   0.2517865006726549   0.5142497089163904   0.6117988035299066   0.13739927331007204   0.8745059205437875   0.13603439643896487   0.024724449844076454   0.6506962545172036   0.9236631370691905   0.727144686907808   0.595813043876427   0.6026640296164473   0.8326616737414118   0.3765538873660493
0.519946486292021   0.9560698219192093   0.5796071033113365   0.8694676560556936   0.07102968335758822   0.9573277381183218   0.22930568623640868   0.617523972451539   0.8780726065068933   0.18394178334860356   0.9775191855637537   0.10327426353514847   0.2662738029769867   0.0465425100385315   0.10301326501996626   0.9672398670961836   0.24154935313291023   0.3958462555213279   0.17935012795077585   0.2400951801883756   0.6457363092564833   0.7931822259048806   0.3466884542093641   0.8635412928223263   0.12578982296446228   0.8371124039856714   0.7670813508980276   0.9940736367666326   0.054760139606874064   0.8797846658673495   0.537775664661619   0.3765496643150937   0.17668753309998078   0.6958428825187459   0.5602564790978652   0.2732754007799452   0.9104137301229941   0.6493003724802144   0.457243214077899   0.30603553368376163   0.6688643769900838   0.2534541169588866   0.27789308612712316   0.06594035349538602   0.023128067733600554   0.4602718910540059   0.931204631917759   0.2023990606730597   0.8973382447691383   0.6231594870683346   0.16412328101973137   0.20832542390642705   0.8425781051622642   0.743374821200985   0.6263476163581124   0.8317757595913333   0.6658905720622834   0.04753193868223902   0.06609113726024714   0.5585003588113882   0.7554768419392893   0.39823156620202455   0.6088479231823481   0.25246482512762647
0.08661246494920552   0.14477744924313796   0.330954837055225   0.18652447163224048   0.06348439721560496   0.6845055581891321   0.39975020513746595   0.9841254109591807   0.16614615244646672   0.06134607112079752   0.2356269241177346   0.7757999870527537   0.3235680472842025   0.3179712499198125   0.6092793077596222   0.9440242274614203   0.6576774752219191   0.27043931123757353   0.5431881704993751   0.38552386865003224   0.9022006332826298   0.872207745035549   0.9343402473170269   0.13305904352240577   0.8155881683334242   0.727430295792411   0.6033854102618019   0.9465345718901653   0.7521037711178192   0.042924737603278966   0.20363520512433592   0.9624091609309845   0.5859576186713525   0.9815786664824815   0.9680082810066013   0.18660917387823084   0.26238957138715   0.663607416562669   0.3587289732469791   0.24258494641681047   0.6047120961652309   0.3931681053250954   0.8155408027476041   0.8570610777667782   0.7025114628826012   0.5209603602895464   0.8812005554305772   0.7240020342443725   0.8869232945491771   0.7935300644971355   0.27781514516877526   0.7774674623542072   0.13481952343135778   0.7506053268938565   0.0741799400444393   0.8150583014232227   0.5488619047600053   0.769026660411375   0.10617165903783797   0.6284491275449918   0.2864723333728552   0.10541924384870609   0.7474426857908588   0.3858641811281813
0.6817602372076242   0.7122511385236107   0.9319018830432548   0.5288031033614031   0.979248774325023   0.19129077823406423   0.05070132761267766   0.8048010691170306   0.09232547977584603   0.39776071373692884   0.7728861824439024   0.027333606762823495   0.9575059563444882   0.6471553868430724   0.6987062423994631   0.21227530533960087   0.408644051584483   0.8781287264316974   0.5925345833616251   0.5838261777946091   0.12217171821162778   0.7727094825829912   0.8450918975707663   0.19796199666642778   0.4404114810040035   0.06045834405938058   0.9131900145275115   0.6691588933050246   0.46116270667898046   0.8691675658253163   0.8624886869148338   0.864357824187994   0.3688372269031344   0.4714068520883875   0.08960250447093143   0.8370242174251705   0.4113312705586462   0.8242514652453151   0.3908962620714683   0.6247489120855696   0.002687218974163194   0.9461227388136179   0.7983616787098431   0.04092273429096054   0.8805155007625354   0.17341325623062656   0.9532697811390768   0.8429607376245328   0.44010401975853186   0.11295491217124598   0.04007976661156529   0.17380184431950813   0.9789413130795515   0.24378734634592963   0.17759107969673144   0.3094440201315141   0.610104086176417   0.7723804942575421   0.08798857522579999   0.4724198027063436   0.19877281561777077   0.948129029012227   0.6970923131543317   0.8476708906207739
0.19608559664360758   0.002006290198609129   0.8987306344444885   0.8067481563298134   0.31557009588107215   0.8285930339679826   0.9454608533054117   0.9637874187052806   0.8754660761225402   0.7156381217967366   0.9053810866938464   0.7899855743857725   0.8965247630429889   0.47185077545080695   0.727790006997115   0.48054155425425843   0.2864206768665719   0.6994702811932648   0.639801431771315   0.008121751547914823   0.08764786124880113   0.7513412521810379   0.9427091186169834   0.16045086092714084   0.8915622646051935   0.7493349619824288   0.043978484172494794   0.3537027045973274   0.5759921687241214   0.9207419280144462   0.09851763086708307   0.38991528589204677   0.700526092601581   0.2051038062177096   0.1931365441732366   0.5999297115062742   0.8040013295585923   0.7332530307669026   0.4653465371761216   0.11938815725201578   0.5175806526920204   0.0337827495736378   0.8255451054048065   0.11126640570410096   0.4299327914432192   0.2824414973925999   0.8828359867878233   0.9508155447769601   0.5383705268380257   0.5331065354101712   0.8388575026153284   0.5971128401796327   0.9623783581139043   0.612364607395725   0.7403398717482453   0.20719755428758593   0.2618522655123232   0.40726080117801533   0.5472033275750088   0.6072678427813117   0.45785093595373094   0.6740077704111127   0.08185679039888714   0.48787968552929595
0.9402702832617106   0.6402250208374749   0.2563116849940806   0.376613279825195   0.5103374918184914   0.35778352344487496   0.37347569820625737   0.4257977350482349   0.9719669649804658   0.8246769880347039   0.5346181955909289   0.8286848948686022   0.009588606866561456   0.21231238063897895   0.7942783238426836   0.6214873405810163   0.7477363413542383   0.8050515794609636   0.24707499626767485   0.01421949779970453   0.28988540540050733   0.13104380904985097   0.16521820586878772   0.5263398122704086   0.3496151221387967   0.49081878821237607   0.9089065208747071   0.14972653244521356   0.8392776303203052   0.1330352647675011   0.5354308226684498   0.7239287973969787   0.8673106653398396   0.30835827673279725   0.0008126270775208003   0.8952439025283764   0.8577220584732781   0.09604589609381829   0.2065343032348372   0.27375656194736014   0.10998571711903982   0.2909943166328547   0.9594593069671624   0.25953706414765565   0.8201003117185325   0.15995050758300372   0.7942411010983746   0.733197251877247   0.47048518957973584   0.6691317193706277   0.8853345802236675   0.5834707194320335   0.6312075592594305   0.5360964546031265   0.3499037575552178   0.8595419220350549   0.763896893919591   0.2277381778703293   0.349091130477697   0.9642980195066785   0.9061748354463129   0.13169228177651102   0.14255682724285978   0.6905414575593183
0.7961891183272731   0.8406979651436564   0.18309752027569742   0.4310043934116627   0.9760888066087406   0.6807474575606526   0.3888564191773228   0.6978071415344156   0.5056036170290048   0.011615738190024998   0.5035218389536552   0.1143364221023821   0.8743960577695743   0.47551928358689843   0.1536180813984374   0.25479450006732723   0.11049916384998325   0.24778110571656917   0.8045269509207404   0.29049648056064875   0.20432432840367032   0.11608882394005815   0.6619701236778807   0.5999550230013304   0.4081352100763972   0.2753908587964018   0.47887260340218324   0.16895062958966778   0.4320464034676566   0.5946434012357492   0.09001618422486045   0.4711434880552522   0.9264427864386517   0.5830276630457242   0.5864943452712053   0.3568070659528701   0.05204672866907752   0.10750837945882571   0.43287626387276784   0.10201256588554286   0.9415475648190943   0.8597272737422565   0.6283493129520273   0.811516085324894   0.737223236415424   0.7436384498021984   0.9663791892741468   0.21156106232356361   0.3290880263390268   0.4682475910057966   0.48750658587196355   0.04261043273389584   0.8970416228713701   0.8736041897700474   0.3974904016471031   0.5714669446786437   0.9705988364327184   0.29057652672432327   0.8109960563758979   0.21465987872577358   0.9185521077636408   0.18306814726549753   0.37811979250313005   0.11264731284023072
0.9770045429445466   0.323340873523241   0.7497704795511027   0.3011312275153366   0.23978130652912263   0.5797024237210425   0.7833912902769559   0.08957016519177301   0.9106932801900959   0.11145483271524598   0.29588470440499237   0.046959732457877164   0.013651657318725703   0.23785064294519856   0.8983943027578892   0.4754927877792335   0.04305282088600731   0.9472741162208753   0.08739824638199144   0.2608329090534599   0.12450071312236644   0.7642059689553777   0.7092784538788615   0.14818559621322921   0.14749617017781982   0.44086509543213676   0.9595079743277588   0.8470543686978925   0.9077148636486972   0.8611626717110942   0.17611668405080289   0.7574842035061196   0.9970215834586014   0.7497078389958483   0.8802319796458106   0.7105244710482425   0.9833699261398756   0.5118571960506497   0.9818376768879212   0.23503168326900892   0.9403171052538684   0.5645830798297744   0.8944394305059299   0.974198774215549   0.8158163921315019   0.8003771108743966   0.18516097662706843   0.8260131780023198   0.668320221953682   0.35951201544225986   0.22565300229930965   0.9789588093044272   0.7606053583049849   0.49834934373116563   0.04953631824850676   0.22147460579830763   0.7635837748463835   0.7486415047353174   0.16930433860269622   0.5109501347500652   0.7802138487065079   0.23678430868466774   0.18746666171477494   0.2759184514810563
0.8398967434526396   0.6722012288548934   0.2930272312088451   0.3017196772655073   0.024080351321137734   0.8718241179804967   0.10786625458177668   0.47570649926318753   0.3557601293674557   0.5123121025382369   0.882213252282467   0.49674768995876034   0.5951547710624708   0.01396275880707129   0.8326769340339603   0.2752730841604527   0.8315709962160873   0.2653212540717539   0.663372595431264   0.7643229494103875   0.05135714750957943   0.028536945387086145   0.4759059337164891   0.4884044979293312   0.21146040405693983   0.35633571653219276   0.18287870250764401   0.18668482066382389   0.1873800527358021   0.484511598551696   0.07501244792586734   0.7109783214006363   0.8316199233683463   0.9721994960134591   0.1927991956434003   0.21423063144187598   0.23646515230587553   0.9582367372063878   0.36012226160944005   0.9389575472814232   0.4048941560897882   0.6929154831346339   0.696749666178176   0.17463459787103575   0.35353700858020876   0.6643785377475477   0.2208437324616869   0.6862300999417045   0.14207660452326892   0.30804282121535503   0.037965029954042884   0.49954527927788067   0.9546965517874668   0.823531222663659   0.9629525820281756   0.7885669578772443   0.12307662841912044   0.8513317266501998   0.7701533863847753   0.5743363264353684   0.8866114761132449   0.893094989443812   0.41003112477533515   0.6353787791539451
0.48171732002345674   0.20017950630917813   0.7132814585971592   0.4607441812829094   0.12818031144324799   0.5358009685616303   0.49243772613547226   0.7745140813412048   0.9861037069199791   0.22775814734627534   0.4544726961814294   0.2749688020633242   0.03140715513251224   0.40422692468261634   0.49152011415325386   0.48640184418607985   0.9083305267133918   0.5528951980324165   0.7213667277684787   0.9120655177507115   0.021719050600146884   0.6598002085886044   0.31133560299314345   0.2766867385967664   0.5400017305766901   0.4596207022794263   0.5980541443959843   0.815942557313857   0.41182141913344217   0.9238197337177959   0.10561641826051202   0.04142847597265219   0.4257177122134631   0.6960615863715206   0.6511437220790827   0.766459673909328   0.39431055708095086   0.29183466168890426   0.15962360792582878   0.2800578297232481   0.48598003036755905   0.7389394636564878   0.43825688015735015   0.3679923119725366   0.46426097976741215   0.07913925506788339   0.12692127716420668   0.09130557337577022   0.924259249190722   0.6195185527884571   0.5288671327682224   0.2753630160619132   0.5124378300572798   0.6956988190706611   0.4232507145077104   0.233934540089261   0.08672011784381677   0.9996372326991405   0.7721069924286278   0.467474866179933   0.692409560762866   0.7078025710102362   0.612483384502799   0.1874170364566849
0.20642953039530687   0.9688631073537485   0.17422650434544887   0.8194247244841483   0.7421685506278948   0.889723852285865   0.04730522718124217   0.728119151108378   0.8179093014371727   0.27020529949740796   0.5184380944130198   0.45275613504646484   0.30547147137989283   0.5745064804267468   0.0951873799053094   0.21882159495720382   0.21875135353607608   0.5748692477276063   0.32308038747668166   0.7513467287772708   0.5263417927732101   0.86706667671737   0.7105970029738826   0.563929692320586   0.31991226237790327   0.8982035693636217   0.5363704986284338   0.7445049678364377   0.5777437117500086   0.008479717077756561   0.48906527144719164   0.01638581672805964   0.7598344103128358   0.7382744175803486   0.9706271770341719   0.5636296816815948   0.454362938932943   0.1637679371536018   0.8754397971288624   0.34480808672439095   0.2356115853968669   0.5888986894259955   0.5523594096521808   0.5934613579471202   0.7092697926236567   0.7218320127086254   0.8417624066782982   0.029531665626534233   0.3893575302457535   0.8236284433450038   0.3053919080498643   0.28502669779009654   0.8116138184957449   0.8151487262672473   0.8163266366026727   0.26864088106203693   0.05177940818290908   0.07687430868689867   0.8456994595685009   0.7050111993804421   0.597416469249966   0.9131063715332969   0.9702596624396385   0.36020311265605115
0.36180488385309917   0.3242076821073014   0.4179002527874576   0.766741754708931   0.6525350912294424   0.6023756693986759   0.5761378461091595   0.7372100890823967   0.2631775609836889   0.7787472260536721   0.2707459380592952   0.4521833912923002   0.45156374248794395   0.9635984997864248   0.45441930145662246   0.18354251023026327   0.3997843343050349   0.8867241910995262   0.6087198418881216   0.47853131084982115   0.8023678650550689   0.9736178195662293   0.6384601794484832   0.11832819819377001   0.44056298120196963   0.6494101374589278   0.2205599266610255   0.35158644348483903   0.7880278899725273   0.047034468060251966   0.644422080551866   0.6143763544024423   0.5248503289888383   0.2682872420065799   0.3736761424925708   0.1621929631101421   0.07328658650089437   0.3046887422201551   0.9192568410359483   0.9786504528798788   0.6735022521958595   0.41796455112062897   0.31053699914782673   0.5001191420300577   0.8711343871407906   0.44434673155439974   0.6720768196993435   0.3817909438362877   0.430571405938821   0.7949365940954719   0.45151689303831805   0.03020450035144867   0.6425435159662938   0.7479021260352199   0.8070948124864521   0.41582814594900636   0.1176931869774554   0.47961488402864   0.43341866999388123   0.25363518283886427   0.04440660047656103   0.1749261418084849   0.5141618289579329   0.27498472995898543
0.37090434828070157   0.756961590687856   0.20362482981010618   0.7748655879289277   0.4997699611399109   0.31261485913345616   0.5315480101107626   0.39307464409264   0.0691985552010899   0.5176782650379843   0.08003111707244455   0.3628701437411913   0.42665503923479614   0.7697761390027644   0.2729363045859925   0.9470419977921849   0.30896185225734074   0.2901612549741245   0.8395176345921113   0.6934068149533207   0.2645552517807797   0.11523511316563957   0.3253558056341783   0.41842208499433525   0.8936509035000781   0.35827352247778366   0.12173097582407214   0.6435564970654075   0.39388094236016724   0.04565866334432747   0.5901829657133095   0.2504818529727676   0.3246823871590774   0.5279803983063431   0.5101518486408649   0.8876117092315763   0.8980273479242812   0.7582042593035787   0.2372155440548725   0.9405697114393913   0.5890654956669404   0.4680430043294542   0.3976979094627613   0.24716289648607065   0.3245102438861607   0.35280789116381467   0.07234210382858296   0.8287408114917354   0.43085934038608253   0.994534368686031   0.9506111280045109   0.18518431442632782   0.03697839802591525   0.9488757053417035   0.3604281622912013   0.9347024614535603   0.7122960108668379   0.4208953070353604   0.8502763136503363   0.047090752221983966   0.8142686629425567   0.6626910477317817   0.6130607695954639   0.10652104078259264
0.22520316727561626   0.19464804340232747   0.21536286013270256   0.859358144296522   0.9006929233894556   0.8418401522385128   0.1430207563041196   0.0306173328047866   0.4698335830033731   0.8473057835524818   0.19240962829960875   0.8454330183784587   0.4328551849774578   0.8984300782107782   0.8319814660084075   0.9107305569248986   0.7205591741106199   0.47753477117541787   0.9817051523580712   0.8636398047029146   0.9062905111680633   0.8148437234436362   0.36864438276260736   0.757118763920322   0.681087343892447   0.6201956800413087   0.1532815226299048   0.8977606196237999   0.7803944205029913   0.7783555278027959   0.010260766325785202   0.8671432868190133   0.3105608374996183   0.9310497442503141   0.8178511380261765   0.02171026844055458   0.8777056525221605   0.03261966603953583   0.985869672017769   0.11097971151565603   0.1571464784115406   0.5550848948641179   0.00416451965969781   0.24733990681274143   0.25085596724347736   0.7402411714204817   0.6355201368970904   0.49022114289241947   0.5697686233510304   0.12004549137917307   0.4822386142671857   0.5924605232686195   0.789374202848039   0.34168996357637715   0.47197784794140046   0.7253172364496061   0.47881336534842067   0.4106402193260631   0.654126709915224   0.7036069680090515   0.6011077128262602   0.37802055328652723   0.668257037897455   0.5926272564933955
0.4439612344147196   0.8229356584224093   0.6640925182377573   0.3452873496806541   0.19310526717124218   0.08269448700192752   0.028572381340666794   0.8550662067882346   0.6233366438202118   0.9626489956227544   0.5463337670734811   0.2626056835196151   0.8339624409721728   0.6209590320463773   0.07435591913208064   0.537288447070009   0.35514907562375203   0.2103188127203142   0.4202292092168566   0.8336814790609575   0.7540413627974919   0.832298259433787   0.7519721713194015   0.24105422256756187   0.3100801283827723   0.009362601011377652   0.08787965308164425   0.8957668728869078   0.11697486121153014   0.9266681140094502   0.05930727174097746   0.04070066609867315   0.49363821739131836   0.9640191183866957   0.5129735046674964   0.7780949825790581   0.6596757764191457   0.3430600863403184   0.4386175855354157   0.24080653550904907   0.30452670079539357   0.13274127362000424   0.018388376318559104   0.40712505644809166   0.5504853379979017   0.30044301418621727   0.2664162049991576   0.1660708338805298   0.2404052096151294   0.2910804131748396   0.17853655191751333   0.27030396099362203   0.12343034840359926   0.3644122991653895   0.11922928017653586   0.22960329489494885   0.6297921310122809   0.4003931807786938   0.6062557755090395   0.45150831231589084   0.9701163545931353   0.05733309443837538   0.1676381899736238   0.21070177680684177
0.6655896537977417   0.9245918208183712   0.1492498136550647   0.80357672035875   0.11510431579983994   0.6241488066321539   0.8828336086559071   0.6375058864782204   0.8746991061847106   0.33306839345731426   0.7042970567383938   0.36720192548459835   0.7512687577811112   0.9686560942919248   0.5850677765618579   0.13759863058964947   0.12147662676883039   0.568262913513231   0.9788120010528184   0.6860903182737587   0.15136027217569514   0.5109298190748556   0.8111738110791946   0.4753885414669169   0.4857706183779535   0.5863379982564845   0.6619239974241299   0.6718118211081667   0.37066630257811356   0.9621891916243306   0.7790903887682228   0.03430593462994645   0.495967196393403   0.6291207981670163   0.07479333202982894   0.6671040091453482   0.7446984386122917   0.6604647038750915   0.489725555467971   0.5295053785556987   0.6232218118434614   0.09220179036186053   0.5109135544151525   0.84341506028194   0.47186153966776617   0.5812719712870049   0.699739743335958   0.36802651881502313   0.9860909212898127   0.9949339730305204   0.0378157459118281   0.6962146977068563   0.6154246187116992   0.032744781406189936   0.25872535714360534   0.6619087630769099   0.11945742231829615   0.40362398323917364   0.18393202511377643   0.9948047539315618   0.3747589837060044   0.7431592793640821   0.6942064696458055   0.46529937537586313
0.7515371718625431   0.6509574890022216   0.18329291523065286   0.6218843150939231   0.2796756321947769   0.06968551771521665   0.4835531718946949   0.2538577962789   0.29358471090496424   0.07475154468469615   0.4457374259828668   0.5576430985720436   0.6781600921932651   0.042006763278506214   0.18701206883926144   0.8957343354951337   0.558702669874969   0.6383827800393326   0.003080043725485017   0.900929581563572   0.1839436861689645   0.8952235006752505   0.3088735740796796   0.43563020618770887   0.4324065143064214   0.24426601167302886   0.1255806588490267   0.8137458910937858   0.15273088211164446   0.1745804939578122   0.6420274869543318   0.5598880948148858   0.8591461712066802   0.09982894927311604   0.196290060971465   0.0022449962428421682   0.18098607901341515   0.05782218599460984   0.00927799213220356   0.10651066074770842   0.6222834091384463   0.4194394059552773   0.006197948406718542   0.20558107918413643   0.4383397229694817   0.5242159052800268   0.697324374327039   0.7699508729964275   0.005933208663060306   0.27994989360699796   0.5717437154780123   0.9562049819026418   0.8532023265514158   0.10536939964918576   0.9297162285236804   0.396316887087756   0.9940561553447356   0.005540450376069718   0.7334261675522155   0.3940718908449138   0.8130700763313204   0.9477182643814599   0.7241481754200119   0.28756123009720536
0.19078666719287424   0.5282788584261826   0.7179502270132934   0.08198015091306894   0.7524469442233925   0.004062953146155792   0.020625852686254387   0.3120292779166414   0.7465137355603323   0.7241130595391578   0.4488821372082421   0.3558242960139996   0.8933114090089164   0.618743659889972   0.5191659086845617   0.9595074089262436   0.8992552536641808   0.6132032095139023   0.7857397411323462   0.5654355180813299   0.08618517733286034   0.6654849451324425   0.06159156571233432   0.27787428798412456   0.8953985101399861   0.13720608670625983   0.34364133869904095   0.1958941370710556   0.14295156591659355   0.13314313356010404   0.32301548601278657   0.8838648591544143   0.3964378303562613   0.4090300740209462   0.8741333488045444   0.5280405631404146   0.5031264213473449   0.7902864141309742   0.35496744011998277   0.5685331542141708   0.6038711676831641   0.17708320461707183   0.5692276989876366   0.0030976361328409713   0.5176859903503038   0.5115982594846293   0.5076361332753022   0.7252233481487165   0.6222874802103177   0.37439217277836956   0.1639947945762613   0.5293292110776608   0.47933591429372413   0.24124903921826552   0.8409793085634747   0.6454643519232466   0.08289808393746283   0.8322189651973193   0.9668459597589303   0.11742378878283204   0.5797716625901179   0.04193255106634511   0.6118785196389475   0.5488906345686612
0.9759004949069539   0.8648493464492732   0.04265082065131091   0.5457929984358202   0.45821450455665   0.3532510869646439   0.5350146873760087   0.8205696502871037   0.8359270243463324   0.9788589141862744   0.37101989279974734   0.2912404392094429   0.3565911100526082   0.7376098749680089   0.5300405842362726   0.6457760872861963   0.27369302611514534   0.9053909097706896   0.5631946244773424   0.5283522985033643   0.6939213635250274   0.8634583587043444   0.9513161048383949   0.9794616639347031   0.7180208686180737   0.9986090122550711   0.908665284187084   0.43366866549888294   0.25980636406142366   0.6453579252904272   0.3736505968110753   0.6130990152117792   0.4238793397150913   0.666499011104153   0.0026307040113279717   0.3218585760023363   0.06728822966248311   0.9288891361361441   0.47259011977505533   0.67608248871614   0.7935952035473377   0.02349822636545454   0.9093954952977129   0.14773019021277564   0.09967384002231028   0.16003986766111009   0.958079390459318   0.1682685262780725   0.3816529714042366   0.1614308554060389   0.04941410627223403   0.7345998607791895   0.12184660734281298   0.5160729301156116   0.6757635094611587   0.12150084556741031   0.6979672676277217   0.8495739190114587   0.6731328054498307   0.799642269565074   0.6306790379652386   0.9206847828753146   0.2005426856747754   0.12355978084893408
0.8370838344179008   0.89718655650986   0.2911471903770625   0.9758295906361585   0.7374099943955905   0.73714668884875   0.33306779991774443   0.807561064358086   0.3557570229913539   0.575715833442711   0.2836536936455104   0.07296120357889642   0.23391041564854095   0.059642903327099414   0.6078901841843517   0.9514603580114861   0.5359431480208193   0.21006898431564072   0.934757378734521   0.15181808844641206   0.9052641100555807   0.2893842014403261   0.7342146930597456   0.028258307597477973   0.06818027563767988   0.39219764493046605   0.44306750268268313   0.05242871696131953   0.33077028124208935   0.6550509560817162   0.10999970276493867   0.2448676526032336   0.9750132582507354   0.07933512263900507   0.8263460091194282   0.17190644902433716   0.7411028426021945   0.019692219311905648   0.21845582493507656   0.22044609101285106   0.2051596945813752   0.8096232349962649   0.28369844620055557   0.06862800256643901   0.29989558452579446   0.5202390335559388   0.54948375314081   0.040369694968961034   0.2317153088881146   0.12804138862547274   0.10641625045812689   0.9879409780076415   0.9009450276460252   0.4729904325437566   0.9964165476931882   0.743073325404408   0.9259317693952899   0.39365530990475156   0.17007053857375995   0.5711668763800708   0.1848289267930954   0.3739630905928459   0.9516147136386834   0.3507207853672197
0.9796692322117202   0.564339855596581   0.6679162674381278   0.28209278280078065   0.6797736476859257   0.04410082204064218   0.11843251429731781   0.24172308783181964   0.4480583387978111   0.9160594334151695   0.012016263839190924   0.25378210982417815   0.5471133111517859   0.4430690008714128   0.015599716146002706   0.5107087844197702   0.621181541756496   0.049413690966661275   0.8455291775722428   0.9395419080396995   0.4363526149634006   0.6754506003738153   0.8939144639335593   0.5888211226724798   0.4566833827516804   0.11111074477723439   0.22599819649543154   0.3067283398716991   0.7769097350657547   0.06700992273659222   0.10756568219811374   0.06500525203987946   0.3288513962679436   0.15095048932142277   0.09554941835892282   0.8112231422157014   0.7817380851161577   0.70788148845001   0.07994970221292011   0.3005143577959311   0.1605565433596617   0.6584677974833486   0.23442052464067736   0.36097244975623166   0.7242039283962611   0.9830171971095333   0.340506060707118   0.7721513270837519   0.2675205456445807   0.8719064523322989   0.11450786421168645   0.4654229872120528   0.490610810578826   0.8048965295957067   0.006942182013572703   0.40041773517217333   0.16175941431088245   0.6539460402742839   0.9113927636546499   0.589194592956472   0.38002132919472476   0.946064551824274   0.8314430614417297   0.28868023516054087
0.21946478583506301   0.28759675434092535   0.5970225368010524   0.9277077854043092   0.49526085743880194   0.3045795572313921   0.2565164760939344   0.1555564583205573   0.22774031179422122   0.43267310489909316   0.142008611882248   0.6901334711085045   0.7371295012153952   0.6277765753033865   0.1350664298686753   0.2897157359363312   0.5753700869045127   0.9738305350291026   0.2236736662140254   0.7005211429798592   0.19534875770978805   0.027765983204828586   0.3922306047722956   0.4118409078193183   0.975883971874725   0.7401692288639032   0.7952080679712432   0.4841331224150091   0.4806231144359231   0.43558967163251117   0.5386915918773088   0.3285766640944518   0.2528828026417019   0.0029165667334180084   0.39668297999506075   0.6384431929859473   0.5157533014263067   0.3751399914300315   0.26161655012638546   0.34872745704961605   0.9403832145217939   0.40130945640092897   0.03794288391236007   0.6482063140697569   0.7450344568120059   0.3735434731961004   0.6457122791400645   0.23636540625043856   0.7691504849372808   0.6333742443321971   0.8505042111688212   0.7522322838354294   0.2885273705013577   0.19778457269968594   0.3118126192915125   0.42365561974097765   0.035644567859655814   0.1948680059662679   0.9151296392964517   0.7852124267550304   0.5198912664333492   0.8197280145362364   0.6535130891700662   0.43648496970541434
0.5795080519115553   0.4184185581353075   0.6155702052577062   0.7882786556356575   0.8344735950995494   0.04487508493920712   0.9698579261176418   0.5519132493852189   0.06532311016226866   0.41150084060701   0.11935371494882048   0.7996809655497894   0.776795739660911   0.21371626790732406   0.807541095657308   0.37602534580881175   0.7411511718012551   0.018848261941056155   0.8924114563608563   0.5908129190537814   0.221259905367906   0.19912024740481976   0.23889836719079   0.15432794934836708   0.6417518534563507   0.7807016892695123   0.6233281619330838   0.3660492937127096   0.8072782583568012   0.7358266043303051   0.6534702358154421   0.8141360443274908   0.7419551481945326   0.32432576372329514   0.5341165208666216   0.0144550787777013   0.9651594085336216   0.11060949581597108   0.7265754252093136   0.6384297329688895   0.22400823673236647   0.09176123387491493   0.8341639688484573   0.047616813915108136   0.002748331364460485   0.8926409864700952   0.5952656016576673   0.8932888645667411   0.3609964779081098   0.1119392972005829   0.9719374397245835   0.5272395708540314   0.5537182195513085   0.3761126928702777   0.31846720390914146   0.7131035265265407   0.811763071356776   0.051786929146982574   0.7843506830425199   0.6986484477488394   0.8466036628231544   0.9411774333310114   0.057775257833206244   0.06021871477994989
0.6225954260907879   0.8494161994560966   0.2236112889847489   0.012601900864841753   0.6198470947263274   0.9567752129860013   0.6283456873270816   0.11931303629810068   0.2588506168182176   0.8448359157854185   0.656408247602498   0.5920734654440692   0.705132397266909   0.46872322291514074   0.33794104369335665   0.8789699389175285   0.8933693259101331   0.41693629376815816   0.5535903606508368   0.18032149116868912   0.04676566308697878   0.47575886043714666   0.4958151028176305   0.12010277638873923   0.42417023699619094   0.6263426609810501   0.2722038138328816   0.10750087552389748   0.8043231422698636   0.6695674479950487   0.6438581265058001   0.9881878392257968   0.5454725254516459   0.8247315322096302   0.987449878903302   0.39611437378172754   0.8403401281847369   0.35600830929448957   0.6495088352099454   0.517144434864199   0.9469708022746038   0.9390720155263313   0.0959184745591086   0.3368229436955099   0.900205139187625   0.46331315508918475   0.6001033717414781   0.21672016730677068   0.47603490219143413   0.8369704941081346   0.32789955790859643   0.10921929178287322   0.6717117599215705   0.16740304611308585   0.6840414314027964   0.12103145255707642   0.12623923446992458   0.34267151390345557   0.6965915524994943   0.7249170787753488   0.28589910628518767   0.986663204608966   0.04708271728954895   0.20777264391114986
0.3389283040105838   0.0475911890826346   0.9511642427304403   0.8709497002156399   0.4387231648229588   0.5842780339934499   0.3510608709889623   0.6542295329088692   0.9626882626315246   0.7473075398853153   0.023161313080365894   0.545010241125996   0.2909765027099541   0.5799044937722294   0.33911988167756957   0.4239787885689196   0.16473726824002952   0.2372329798687739   0.6425283291780752   0.6990617097935707   0.8788381619548419   0.2505697752598079   0.5954456118885263   0.4912890658824209   0.539909857944258   0.2029785861771733   0.6442813691580859   0.6203393656667809   0.10118669312129926   0.6187005521837234   0.2932204981691236   0.9661098327579117   0.1384984304897746   0.8713930122984082   0.2700591850887577   0.4210995916319157   0.8475219277798205   0.2914885185261787   0.9309393034111881   0.9971208030629961   0.682784659539791   0.054255538657404796   0.28841097423311296   0.29805909326942537   0.8039464975849491   0.8036857633975969   0.6929653623445867   0.8067700273870045   0.264036639640691   0.6007071772204237   0.04868399318650076   0.1864306617202236   0.16284994651939178   0.9820066250367002   0.7554634950173772   0.2203208289623119   0.024351516029617177   0.11061361273829207   0.48540430992861944   0.7992212373303962   0.1768295882497967   0.8191250942121133   0.5544650065174312   0.8021004342674001
0.4940449287100057   0.7648695555547086   0.26605403228431834   0.5040413409979747   0.6900984311250566   0.9611837921571117   0.5730886699397316   0.6972713136109702   0.4260617914843656   0.3604766149366881   0.5244046767532309   0.5108406518907466   0.26321184496497385   0.37846998989998787   0.7689411817358538   0.2905198229284347   0.23886032893535666   0.2678563771616958   0.2835368718072343   0.4912985855980385   0.06203074068555998   0.4487312829495824   0.7290718652898031   0.6891981513306384   0.5679858119755542   0.6838617273948738   0.4630178330054847   0.18515681033266368   0.8778873808504976   0.7226779352377621   0.889929163065753   0.48788549672169346   0.451825589366132   0.3622013203010741   0.36552448631252216   0.9770448448309469   0.18861374440115813   0.9837313304010862   0.5965833045766684   0.6865250219025122   0.9497534154658015   0.7158749532393904   0.31304643276943406   0.19522643630447364   0.8877226747802415   0.26714367028980796   0.5839745674796311   0.5060282849738352   0.3197368628046872   0.5832819428949341   0.12095673447414636   0.32087147464117155   0.44184948195418966   0.8606040076571719   0.23102757140839333   0.832985977919478   0.9900238925880577   0.49840268735609783   0.8655030850958711   0.8559411330885313   0.8014101481868996   0.5146713569550116   0.2689197805192028   0.16941611118601904
0.8516567327210981   0.7987964037156212   0.9558733477497687   0.9741896748815454   0.9639340579408566   0.5316527334258133   0.3718987802701377   0.46816138990771017   0.6441971951361694   0.9483707905308791   0.25094204579599133   0.1472899152665386   0.20234771318197972   0.08776678287370723   0.019914474387598004   0.3143039373470605   0.21232382059392205   0.5893640955176094   0.15441138929172682   0.45836280425852927   0.4109136724070225   0.07469273856259777   0.885491608772524   0.28894669307251025   0.5592569396859244   0.2758963348469765   0.9296182610227552   0.31475701819096485   0.5953228817450678   0.7442436014211633   0.5577194807526176   0.8465956282832547   0.9511256866088984   0.795872810890284   0.3067774349566263   0.6993057130167161   0.7487779734269187   0.7081060280165768   0.28686296056902827   0.3850017756696556   0.5364541528329967   0.11874193249896745   0.13245157127730145   0.9266389714111263   0.12554048042597415   0.044049193936369684   0.24695996250477745   0.6376922783386161   0.5662835407400497   0.7681528590893931   0.3173417014820222   0.3229352601476512   0.970960658994982   0.02390925766822989   0.7596222207294046   0.47633963186439654   0.01983497238608351   0.2280364467779458   0.4528447857727783   0.7770339188476805   0.2710569989591648   0.5199304187613689   0.16598182520375004   0.3920321431780248
0.7346028461261681   0.4011884862624015   0.03353025392644858   0.46539317176689854   0.609062365700194   0.3571392923260318   0.7865702914216711   0.8277008934282825   0.042778824960144256   0.5889864332366387   0.46922858993964894   0.5047656332806312   0.07181816596516231   0.5650771755684088   0.7096063692102444   0.028426001416234668   0.0519831935790788   0.337040728790463   0.2567615834374661   0.2513920825685542   0.780926194619914   0.8171103100290941   0.09077975823371606   0.8593599393905293   0.04632334849374584   0.4159218237666925   0.05724950430726748   0.39396676762363086   0.43726098279355186   0.05878253144066068   0.2706792128855963   0.5662658741953485   0.39448215783340757   0.469796098204022   0.8014506229459474   0.06150024091471723   0.3226639918682453   0.9047189226356132   0.09184425373570297   0.03307423949848256   0.27068079828916647   0.5676781938451503   0.8350826702982369   0.7816821569299284   0.48975460366925244   0.7505678838160562   0.7443029120645208   0.9223222175393989   0.44343125517550663   0.3346460600493637   0.6870534077572533   0.528355449915768   0.006170272381954781   0.275863528608703   0.416374194871657   0.9620895757204196   0.6116881145485472   0.806067430404681   0.6149235719257096   0.9005893348057024   0.2890241226803019   0.9013485077690678   0.5230793181900066   0.8675150953072198
0.018343324391135472   0.3336703139239176   0.6879966478917697   0.0858329383772915   0.528588720721883   0.5831024301078613   0.9436937358272489   0.16351072083789256   0.08515746554637639   0.2484563700584977   0.2566403280699956   0.6351552709221245   0.0789871931644216   0.9725928414497946   0.8402661331983386   0.6730656952017049   0.4672990786158744   0.16652541104511362   0.22534256127262903   0.7724763603960025   0.17827495593557247   0.2651769032760458   0.7022632430826224   0.9049612650887827   0.159931631544437   0.9315065893521282   0.01426659519085266   0.8191283267114912   0.631342910822554   0.3484041592442668   0.07057285936360372   0.6556176058735986   0.5461854452761776   0.09994778918576915   0.8139325312936081   0.020462334951474127   0.467198252111756   0.1273549477359745   0.9736663980952694   0.3473966397497692   0.9998991734958816   0.9608295366908609   0.7483238368226405   0.5749202793537667   0.8216242175603091   0.6956526334148151   0.04606059374001803   0.6699590142649839   0.6616925860158721   0.7641460440626868   0.03179399854916536   0.8508306875534928   0.030349675193318132   0.41574188481842006   0.9612211391855616   0.19521308167989412   0.48416422991714053   0.3157940956326509   0.14728860789195353   0.17475074672841998   0.016965977805384527   0.1884391478966764   0.17362220979668408   0.8273541069786507
0.017066804309502935   0.22760961120581552   0.4252983729740436   0.2524338276248841   0.19544258674919382   0.5319569777910005   0.37923777923402563   0.5824748133599001   0.5337500007333217   0.7678109337283135   0.34744378068486026   0.7316441258064074   0.5034003255400036   0.35206904890989354   0.3862226414992986   0.5364310441265132   0.019236095622863037   0.03627495327724264   0.23893403360734505   0.36168029739809326   0.0022701178174785097   0.8478358053805662   0.06531182381066099   0.5343261904194425   0.9852033135079755   0.6202261941747508   0.6400134508366173   0.28189236279455837   0.7897607267587817   0.0882692163837503   0.26077567160259174   0.6994175494346583   0.25601072602546004   0.32045828265543674   0.9133318909177315   0.9677734236282509   0.7526104004854565   0.9683892337455432   0.527109249418433   0.43134237950173765   0.7333743048625935   0.9321142804683006   0.28817521581108785   0.06966208210364441   0.7311041870451149   0.08427847508773433   0.22286339200042687   0.5353358916842019   0.7459008735371394   0.4640522809129836   0.5828499411638095   0.25344352888964355   0.9561401467783576   0.37578306452923327   0.32207426956121776   0.5540259794549852   0.7001294207528975   0.055324781873796545   0.4087423786434862   0.5862525558267343   0.9475190202674411   0.08693554812825333   0.8816331292250533   0.15491017632499668
0.21414471540484759   0.15482126765995274   0.5934579134139655   0.08524809422135227   0.48304052835973266   0.07054279257221842   0.3705945214135386   0.5499122025371503   0.7371396548225932   0.6064905116592348   0.787744580249729   0.29646867364750684   0.7809995080442357   0.23070744713000155   0.4656703106885113   0.7424426941925215   0.08087008729133809   0.175382665256205   0.05692793204502505   0.1561901383657872   0.13335106702389704   0.08844711712795167   0.17529480281997173   0.0012799620407905397   0.9192063516190494   0.933625849467999   0.5818368894060063   0.9160318678194382   0.4361658232593168   0.8630830568957805   0.21124236799246768   0.3661196652822879   0.6990261684367235   0.2565925452365457   0.4234977877427386   0.0696509916347811   0.9180266603924879   0.025885098106544137   0.9578274770542273   0.32720829744225954   0.8371565731011498   0.8505024328503391   0.9008995450092022   0.1710181590764723   0.7038055060772528   0.7620553157223875   0.7256047421892305   0.16973819703568177   0.7845991544582033   0.8284294662543885   0.1437678527832243   0.25370632921624353   0.34843333119888653   0.965346409358608   0.9325254847907566   0.8875866639339556   0.649407162762163   0.7087538641220623   0.509027697048018   0.8179356722991745   0.7313805023696751   0.6828687660155182   0.5512002199937907   0.490727374856915
0.8942239292685252   0.832366333165179   0.6503006749845884   0.31970921578044265   0.1904184231912725   0.07031101744279161   0.9246959327953579   0.14997101874476088   0.40581926873306917   0.24188155118840307   0.7809280800121335   0.8962646895285173   0.05738593753418267   0.27653514182979505   0.848402595221377   0.008678025594561775   0.40797877477201966   0.5677812777077327   0.3393748981733589   0.19074235329538727   0.6765982724023446   0.8849125116922145   0.7881746781795682   0.7000149784384723   0.7823743431338193   0.05254617852703541   0.13787400319497986   0.3803057626580297   0.5919559199425468   0.9822351610842438   0.213178070399622   0.2303347439132688   0.18613665120947762   0.7403536098958408   0.43224999038748846   0.33407005438475146   0.12875071367529495   0.46381846806604565   0.5838473951661115   0.32539202879018964   0.7207719389032753   0.896037190358313   0.24447249699275253   0.1346496754948024   0.04417366650093066   0.011124678666098477   0.45629781881318426   0.43463469705633007   0.26179932336711137   0.9585785001390631   0.31842381561820443   0.05432893439830038   0.6698434034245645   0.9763433390548193   0.10524574521858243   0.8239941904850315   0.4837067522150869   0.23598972915897856   0.672995754831094   0.4899241361002801   0.35495603853979196   0.7721712610929329   0.08914835966498251   0.1645321073100905
0.6341840996365168   0.8761340707346199   0.8446758626722299   0.029882431815288105   0.5900104331355861   0.8650093920685215   0.3883780438590457   0.5952477347589581   0.32821110976847473   0.9064308919294584   0.06995422824084126   0.5409188003606576   0.6583677063439102   0.9300875528746391   0.9647084830222589   0.7169246098756261   0.17466095412882326   0.6940978237156605   0.29171272819116484   0.22700047377534593   0.8197049155890312   0.9219265626227277   0.20256436852618231   0.06246836646525546   0.18552081595251455   0.04579249188810771   0.3578885058539524   0.032585934649967355   0.5955103828169285   0.18078309981958623   0.9695104619949066   0.4373381998910093   0.26729927304845374   0.2743522078901279   0.8995562337540655   0.8964193995303517   0.6089315667045435   0.34426465501548875   0.9348477507318066   0.17949478965472557   0.4342706125757203   0.6501668312998282   0.6431350225406418   0.9524943158793796   0.6145656969866891   0.7282402686771006   0.44057065401445944   0.8900259494141242   0.4290448810341745   0.6824477767889928   0.08268214816050708   0.8574400147641568   0.833534498217246   0.5016646769694065   0.1131716861656004   0.4201018148731475   0.5662352251687923   0.2273124690792787   0.21361545241153498   0.5236824153427958   0.9573036584642487   0.88304781406379   0.27876770167972836   0.3441876256880703
0.5230330458885285   0.23288098276396182   0.6356326791390866   0.39169330980869066   0.9084673489018394   0.5046407140868613   0.19506202512462717   0.5016673603945665   0.47942246786766496   0.8221929372978685   0.11237987696412009   0.6442273456304097   0.645887969650419   0.3205282603284619   0.9992081907985197   0.22412553075726224   0.07965274448162671   0.09321579124918317   0.7855927383869847   0.7004431154144664   0.12234908601737797   0.21016797718539318   0.5068250367072563   0.3562554897263961   0.5993160401288495   0.9772869944214314   0.8711923575681697   0.9645621799177054   0.6908486912270101   0.47264628033457007   0.6761303324435426   0.4628948195231389   0.21142622335934508   0.6504533430367017   0.5637504554794225   0.8186674738927292   0.5655382537089261   0.3299250827082397   0.5645422646809027   0.5945419431354669   0.4858855092272994   0.23670929145905656   0.7789495262939181   0.8940988277210006   0.3635364232099214   0.026541314273663404   0.27212448958666174   0.5378433379946045   0.7642203830810719   0.04925431985223205   0.400932132018492   0.5732811580768991   0.07337169185406185   0.5766080395176619   0.7248017995749494   0.11038633855376015   0.8619454684947168   0.9261546964809604   0.16105134409552696   0.291718864661031   0.2964072147857907   0.5962296137727207   0.5965090794146242   0.6971769215255641
0.8105217055584912   0.35952032231366404   0.817559553120706   0.8030780938045635   0.4469852823485699   0.33297900804000063   0.5454350635340444   0.2652347558099591   0.682764899267498   0.2837246881877686   0.1445029315155524   0.6919535977330601   0.609393207413436   0.7071166486701066   0.419701131940603   0.5815672591792999   0.7474477389187193   0.7809619521891463   0.25864978784507603   0.2898483945182689   0.45104052413292867   0.18473233841642564   0.6621407084304518   0.5926714729927048   0.6405188185744374   0.8252120161027616   0.8445811553097458   0.7895933791881413   0.19353353622586753   0.49223300806276093   0.29914609177570134   0.5243586233781823   0.5107686369583696   0.20850831987499233   0.15464316026014896   0.8324050256451222   0.9013754295449334   0.5013916712048857   0.734942028319546   0.25083776646582234   0.15392769062621417   0.7204297190157395   0.47629224047447   0.9609893719475534   0.7028871664932855   0.5356973805993138   0.8141515320440181   0.36831789895484857   0.06236834791884814   0.7104853644965522   0.9695703767342724   0.5787245197667072   0.8688348116929806   0.21825235643379126   0.670424284958571   0.05436589638852501   0.35806617473461105   0.009744036558798918   0.5157811246984221   0.22196087074340282   0.45669074518967756   0.5083523653539133   0.780839096378876   0.9711231042775805
0.3027630545634634   0.7879226463381738   0.30454685590440606   0.010133732330027078   0.5998758880701779   0.25222526573886   0.4903953238603879   0.6418158333751786   0.5375075401513297   0.5417399012423078   0.5208249471261156   0.06309131360847126   0.6686727284583491   0.32348754480851655   0.8504006621675446   0.00872541721994624   0.3106065537237381   0.31374350824971764   0.33461953746912254   0.7867645464765435   0.8539158085340606   0.8053911428958044   0.5537804410902465   0.815641442198963   0.5511527539705972   0.017468496557630633   0.24923358518584046   0.8055077098689358   0.9512768659004193   0.7652432308187707   0.7588382613254525   0.16369187649375735   0.4137693257490895   0.22350332957646285   0.23801331419933694   0.10060056288528611   0.7450965972907404   0.9000157847679463   0.38761265203179235   0.09187514566533987   0.43449004356700227   0.5862722765182287   0.0529931145626698   0.30511059918879646   0.5805742350329417   0.7808811336224243   0.49921267347242326   0.4894691569898335   0.029421481062344625   0.7634126370647937   0.24997908828658283   0.6839614471208977   0.07814461516192539   0.998169406246023   0.4911408269611303   0.5202695706271403   0.6643752894128359   0.7746660766695601   0.25312751276179335   0.41966900774185417   0.9192786921220956   0.8746502919016138   0.8655148607300011   0.3277938620765143
0.4847886485550933   0.28837801538338514   0.8125217461673312   0.02268326288771785   0.9042144135221515   0.5074968817609609   0.31330907269490793   0.5332141058978843   0.8747929324598069   0.7440842446961672   0.06332998440832512   0.8492526587769867   0.7966483172978815   0.7459148384501442   0.5721891574471948   0.32898308814984645   0.1322730278850456   0.971248761780584   0.31906164468540144   0.9093140804079923   0.21299433576295007   0.09659846987897015   0.4535467839554004   0.581520218331478   0.7282056872078568   0.808220454495585   0.6410250377880692   0.5588369554437602   0.8239912736857052   0.30072357273462413   0.32771596509316125   0.025622849545875813   0.9491983412258984   0.556639328038457   0.26438598068483615   0.17637019076888907   0.15255002392801686   0.8107244895883128   0.6921968232376413   0.8473871026190426   0.02027699604297125   0.8394757278077288   0.37313517855223993   0.9380730222110504   0.8072826602800212   0.7428772579287587   0.9195883945968395   0.35655280387957233   0.0790769730721644   0.9346568034331737   0.2785633568087703   0.7977158484358121   0.25508569938645914   0.6339332306985495   0.9508473917156091   0.7720929988899363   0.30588735816056073   0.07729390266009252   0.686461411030773   0.5957228081210473   0.1533373342325439   0.2665694130717797   0.9942645877931316   0.7483357055020046
0.13306033818957264   0.4270936852640509   0.6211294092408917   0.8102626832909543   0.3257776779095515   0.6842164273352922   0.7015410146440522   0.45370987941138197   0.24670070483738707   0.7495596239021186   0.42297765783528185   0.6559940309755699   0.991615005450928   0.11562639320356906   0.4721302661196728   0.8839010320856335   0.6857276472903672   0.03833249054347654   0.7856688550888998   0.28817822396458626   0.5323903130578233   0.7717630774716968   0.7914042672957683   0.5398425184625817   0.39932997486825067   0.3446693922076459   0.1702748580548766   0.7295798351716274   0.0735522969586992   0.6604529648723537   0.4687338434108244   0.27586995576024537   0.8268515921213121   0.9108933409702351   0.045756185575542535   0.6198759247846756   0.8352365866703843   0.7952669477666661   0.5736259194558697   0.735974892699042   0.14950893938001703   0.7569344572231895   0.7879570643669699   0.4477966687344558   0.6171186263221937   0.9851713797514927   0.9965527970712016   0.9079541502718741   0.21778865145394305   0.6405019875438468   0.826277939016325   0.17837431510024673   0.14423635449524386   0.9800490226714931   0.3575440956055006   0.9025043593400013   0.3173847623739317   0.06915568170125791   0.31178791002995804   0.28262843455532577   0.4821481757035475   0.2738887339345918   0.7381619905740883   0.5466535418562838
0.3326392363235305   0.5169542767114023   0.9502049262071185   0.09885687312182798   0.7155206100013368   0.5317828969599095   0.9536521291359169   0.19090272284995388   0.4977319585473937   0.8912809094160627   0.1273741901195919   0.012528407749707163   0.35349560405214986   0.9112318867445697   0.7698300945140913   0.11002404840970584   0.036110841678218174   0.8420762050433118   0.45804218448413325   0.8273956138543801   0.5539626659746707   0.5681874711087199   0.719880193910045   0.2807420719980963   0.22132342965114019   0.051233194397317695   0.7696752677029265   0.18188519887626833   0.5058028196498034   0.5194502974374081   0.8160231385670097   0.9909824760263144   0.008070861102409673   0.6281693880213455   0.6886489484474178   0.9784540682766073   0.6545752570502598   0.7169375012767757   0.9188188539333265   0.8684300198669015   0.6184644153720417   0.874861296233464   0.4607766694491932   0.041034406012521396   0.06450174939737095   0.306673825124744   0.7408964755391482   0.7602923340144251   0.8431783197462308   0.25544063072742634   0.9712212078362217   0.5784071351381568   0.33737550009642736   0.7359903332900182   0.15519806926921204   0.5874246591118423   0.3293046389940177   0.10782094526867274   0.4665491208217942   0.6089705908352351   0.6747293819437579   0.390883443991897   0.5477302668884678   0.7405405709683336
0.056264966571716285   0.516022147758433   0.08695359743927458   0.6995061649558122   0.9917632171743453   0.209348322633689   0.3460571219001264   0.9392138309413871   0.14858489742811454   0.9539076919062627   0.37483591406390465   0.3608066958032303   0.8112093973316872   0.2179173586162445   0.21963784479469264   0.773382036691388   0.48190475833766944   0.11009641334757178   0.7530887239728984   0.164411445856153   0.8071753763939116   0.7192129693556748   0.2053584570844306   0.42387087488781944   0.7509104098221953   0.20319082159724178   0.11840485964515603   0.7243647099320072   0.7591471926478499   0.9938424989635528   0.7723477377450296   0.7851508789906201   0.6105622952197354   0.039934807057290106   0.397511823681125   0.42434418318738976   0.7993528978880482   0.8220174484410456   0.17787397888643236   0.6509621464960017   0.31744813955037876   0.7119210350934738   0.42478525491353397   0.48655070063984873   0.5102727631564672   0.992708065737799   0.21942679782910338   0.06267982575202931   0.7593623533342719   0.7895172441405572   0.10102193818394735   0.3383151158200221   0.00021516068642200349   0.7956747451770045   0.3286742004389177   0.553164236829402   0.3896528654666866   0.7557399381197144   0.9311623767577927   0.12882005364201224   0.5902999675786385   0.9337224896786688   0.7532883978713604   0.4778579071460105
0.27285182802825964   0.22180145458519498   0.32850314295782634   0.9913072065061618   0.7625790648717924   0.22909338884739594   0.10907634512872297   0.9286273807541325   0.0032167115375205   0.4395761447068387   0.008054406944775612   0.5903122649341104   0.0030015508510984968   0.6439013995298342   0.679380206505858   0.0371480281047084   0.6133486853844119   0.8881614614101198   0.7482178297480653   0.9083279744626962   0.02304871780577348   0.954438971731451   0.9949294318767049   0.43047006731668563   0.7501968897775139   0.732637517146256   0.6664262889188786   0.43916286081052386   0.9876178249057214   0.5035441282988601   0.5573499437901557   0.5105354800563914   0.9844011133682009   0.06396798359202141   0.54929553684538   0.920223215122281   0.9813995625171024   0.4200665840621872   0.8699153303395221   0.8830751870175726   0.3680508771326905   0.5319051226520674   0.12169750059145684   0.9747472125548764   0.345002159326917   0.5774661509206164   0.1267680687147519   0.5442771452381907   0.5948052695494032   0.8448286337743603   0.4603417797958733   0.10511428442766689   0.6071874446436818   0.34128450547550027   0.9029918360057176   0.5945788043712755   0.6227863312754809   0.2773165218834789   0.3536962991603377   0.6743555892489945   0.6413867687583785   0.8572499378212917   0.48378096882081556   0.7912804022314219
0.273335891625688   0.32534481516922426   0.3620834682293587   0.8165331896765455   0.9283337322987709   0.7478786642486078   0.2353153995146068   0.27225604443835477   0.33352846274936776   0.9030500304742475   0.7749736197187335   0.1671417600106879   0.726341018105686   0.5617655249987472   0.8719817837130158   0.5725629556394124   0.10355468683020504   0.2844490031152684   0.5182854845526781   0.8982073663904179   0.4621679180718265   0.4271990652939767   0.03450451573186255   0.10692696415899591   0.18883202644613853   0.10185425012475248   0.6724210475025039   0.2903937744824504   0.2604982941473676   0.35397558587614464   0.437105647987897   0.0181377300440956   0.9269698313979998   0.4509255554018971   0.6621320282691635   0.8509959700334077   0.20062881329231386   0.88916003040315   0.7901502445561477   0.2784330143939953   0.09707412646210882   0.6047110272878815   0.27186476000346954   0.38022564800357744   0.6349062083902823   0.17751196199390482   0.237360244271607   0.27329868384458156   0.4460741819441438   0.07565771186915234   0.5649391967691032   0.9829049093621312   0.18557588779677622   0.7216821259930077   0.1278335487812062   0.9647671793180356   0.25860605639877643   0.2707565705911106   0.4657015205120427   0.11377120928462786   0.05797724310646257   0.3815965401879607   0.675551275955895   0.8353381948906325
0.9609031166443538   0.7768855129000791   0.40368651595242544   0.4551125468870551   0.32599690825407146   0.5993735509061744   0.16632627168081843   0.18181386304247352   0.8799227263099276   0.523715839037022   0.6013870749117153   0.19890895368034237   0.6943468385131514   0.8020337130440143   0.47355352613050905   0.2341417743623068   0.435740782114375   0.5312771424529037   0.007852005618466325   0.12037056507767893   0.37776353900791243   0.14968060226494304   0.33230072966257135   0.2850323701870464   0.4168604223635587   0.3727950893648639   0.9286142137101459   0.8299198232999914   0.09086351410948723   0.7734215384586896   0.7622879420293275   0.6481059602575178   0.21094078779955958   0.24970569942166754   0.16090086711761223   0.44919700657717543   0.5165939492864081   0.4476719863776532   0.6873473409871033   0.21505523221486864   0.08085316717203313   0.9163948439247495   0.6794953353686369   0.0946846671371897   0.7030896281641207   0.7667142416598065   0.3471946057060656   0.8096522969501433   0.28622920580056205   0.39391915229494257   0.4185803919959197   0.979732473650152   0.1953656916910748   0.620497613836253   0.6562924499665922   0.3316265133926342   0.9844249038915153   0.3707919144145855   0.49539158284898   0.8824295068154587   0.4678309546051071   0.9231199280369323   0.8080442418618767   0.6673742746005902
0.386977787433074   0.006725084112182775   0.12854890649323988   0.5726896074634005   0.6838881592689533   0.24001084245237633   0.7813543007871743   0.7630373105132572   0.39765895346839125   0.8460916901574338   0.36277390879125465   0.7833048368631051   0.20229326177731644   0.22559407632118073   0.7064814588246624   0.45167832347047093   0.2178683578858012   0.8548021619065952   0.21108987597568243   0.5692488166550121   0.7500374032806941   0.931682233869663   0.4030456341138057   0.901874542054422   0.36305961584762014   0.9249571497574802   0.2744967276205658   0.32918493459102155   0.679171456578667   0.6849463073051039   0.4931424268333915   0.5661476240777644   0.28151250311027565   0.8388546171476701   0.13036851804213684   0.7828427872146593   0.07921924133295924   0.6132605408264894   0.42388705921747444   0.3311644637441884   0.861350883447158   0.7584583789198941   0.21279718324179198   0.7619156470891763   0.11131348016646392   0.8267761450502312   0.8097515491279863   0.8600411050347542   0.7482538643188438   0.901818995292751   0.5352548215074205   0.5308561704437327   0.06908240774017686   0.2168726879876471   0.04211239467402902   0.9647085463659683   0.7875699046299012   0.378018070839977   0.9117438766318922   0.18186575915130893   0.708350663296942   0.7647575300134877   0.4878568174144178   0.8507012954071206
0.8469997798497839   0.006299151093593481   0.27505963417262574   0.08878564831794432   0.73568629968332   0.1795230060433623   0.46530808504463944   0.2287445432831901   0.9874324353644762   0.2777040107506113   0.930053263537219   0.6978883728394575   0.9183500276242994   0.0608313227629642   0.8879408688631899   0.7331798264734892   0.13078012299439817   0.6828132519229871   0.9761969922312977   0.5513140673221802   0.4224294596974562   0.9180557219094996   0.48834017481688   0.7006127719150598   0.5754296798476723   0.9117565708159061   0.21328054064425425   0.6118271235971154   0.8397433801643523   0.7322335647725438   0.7479724555996148   0.38308258031392534   0.8523109447998761   0.45452955402193246   0.8179191920623958   0.6851942074744679   0.9339609171755767   0.39369823125896825   0.9299783231992059   0.9520143810009787   0.8031807941811785   0.710884979335981   0.9537813309679081   0.4007003136787984   0.3807513344837223   0.7928292574264815   0.46544115615102805   0.7000875417637387   0.80532165463605   0.8810726866105755   0.2521606155067738   0.08826041816662328   0.9655782744716976   0.14883912183803163   0.504188159907159   0.7051778378526979   0.1132673296718216   0.6943095678160992   0.6862689678447632   0.019983630378230078   0.17930641249624488   0.3006113365571309   0.7562906446455573   0.06796924937725139
0.37612561831506636   0.5897263572211499   0.8025093136776492   0.667268935698453   0.9953742838313441   0.7968970997946683   0.33706815752662117   0.9671813939347144   0.19005262919529406   0.9158244131840929   0.08490754201984735   0.878920975768091   0.22447435472359636   0.7669852913460613   0.5807193821126884   0.1737431379153931   0.11120702505177477   0.07267572352996209   0.8944504142679252   0.153759507537163   0.9319006125555299   0.7720643869728312   0.1381597696223678   0.08579025815991159   0.5557749942404635   0.18233802975168134   0.3356504559447186   0.4185213224614586   0.5604007104091194   0.385440929957013   0.9985822984180974   0.4513399285267443   0.3703480812138254   0.46961651677292016   0.91367475639825   0.5724189527586533   0.14587372649022906   0.7026312254268589   0.3329553742855617   0.3986758148432602   0.0346667014384543   0.6299555018968968   0.4385049600176366   0.24491630730609718   0.10276608888292443   0.8578911149240657   0.3003451903952688   0.15912604914618558   0.5469910946424609   0.6755530851723842   0.9646947344505502   0.740604726684727   0.9865903842333414   0.29011215521537126   0.9661124360324528   0.28926479815798267   0.616242303019516   0.8204956384424511   0.052437679634202775   0.7168458453993294   0.47036857652928693   0.11786441301559221   0.719482305348641   0.31817003055606924
0.43570187509083264   0.4879089111186954   0.28097734533100444   0.07325372324997206   0.33293578620790826   0.6300177961946298   0.9806321549357356   0.9141276741037865   0.7859446915654473   0.9544647110222455   0.015937420485185386   0.1735229474190595   0.7993543073321059   0.6643525558068742   0.049824984452732556   0.8842581492610768   0.18311200431258987   0.8438569173644231   0.9973873048185298   0.16741230386174735   0.7127434277833029   0.725992504348831   0.2779049994698887   0.8492422733056781   0.27704155269247027   0.2380835932301356   0.9969276541388843   0.775988550055706   0.944105766484562   0.6080657970355058   0.016295499203148673   0.8618608759519196   0.15816107491911469   0.6536010860132603   0.00035807871796328774   0.6883379285328601   0.3588067675870088   0.989248530206386   0.9505330942652307   0.8040797792717833   0.17569476327441896   0.1453916128419628   0.9531457894467009   0.6366674754100359   0.46295133549111606   0.41939910849313183   0.6752407899768123   0.7874252021043578   0.18590978279864578   0.18131551526299625   0.678313135837928   0.011436652048651763   0.24180401631408377   0.5732497182274905   0.6620176366347792   0.1495757760967322   0.08364294139496907   0.9196486322142302   0.661659557916816   0.4612378475638721   0.7248361738079603   0.9304001020078442   0.7111264636515853   0.6571580682920888
0.5491414105335413   0.7850084891658814   0.7579806742048842   0.020490592882052894   0.08619007504242526   0.3656093806727495   0.08273988422807205   0.2330653907776951   0.9002802922437795   0.1842938654097533   0.40442674839014414   0.22162873872904332   0.6584762759296957   0.6110441471822629   0.7424091117553648   0.07205296263231113   0.5748333345347266   0.6913955149680326   0.08074955383854893   0.610815115068439   0.8499971607267663   0.7609954129601886   0.3696230901869637   0.9536570467763502   0.3008557501932251   0.9759869237943072   0.6116424159820795   0.9331664538942973   0.2146656751507998   0.6103775431215577   0.5289025317540074   0.7001010631166023   0.31438538290702034   0.42608367771180433   0.12447578336386327   0.47847232438755893   0.6559091069773246   0.8150395305295415   0.3820666716084984   0.4064193617552478   0.08107577244259799   0.12364401556150884   0.30131711776994946   0.7956042466868087   0.23107861171583163   0.3626486026013203   0.9316940275829857   0.8419471999104585   0.9302228615226066   0.38666167880701313   0.3200516116009063   0.9087807460161612   0.7155571863718068   0.7762841356854555   0.7911490798468989   0.20867968289955902   0.4011718034647865   0.3502004579736511   0.6666732964830356   0.7302073585120001   0.7452626964874619   0.5351609274441096   0.28460662487453725   0.3237879967567523
0.6641869240448639   0.41151691188260076   0.9832895071045878   0.5281837500699436   0.43310831232903224   0.04886830928128048   0.05159547952160205   0.686236550159485   0.5028854508064257   0.6622066304742673   0.7315438679206957   0.7774558041433237   0.7873282644346189   0.8859224947888119   0.9403947880737968   0.5687761212437648   0.38615646096983236   0.5357220368151607   0.27372149159076126   0.8385687627317646   0.6408937644823706   0.0005611093710511331   0.989114866716224   0.5147807659750123   0.9767068404375067   0.5890441974884504   0.005825359611636204   0.9865970159050688   0.5435985281084744   0.5401758882071699   0.9542298800900342   0.3003604657455837   0.04071307730204876   0.8779692577329026   0.2226860121693384   0.52290466160226   0.2533848128674299   0.9920467629440907   0.2822912240955415   0.9541285403584953   0.8672283518975975   0.4563247261289299   0.008569732504780301   0.11555977762673066   0.22633458741522702   0.4557636167578788   0.019454865788556305   0.6007790116517183   0.2496277469777204   0.8667194192694284   0.013629506176920101   0.6141819957466496   0.706029218869246   0.32654353106225853   0.05939962608688595   0.3138215300010659   0.6653161415671972   0.448574273329356   0.8367136139175475   0.7909168683988058   0.4119313286997673   0.4565275103852654   0.554422389822006   0.8367883280403106
0.5447029768021697   0.00020278425633547164   0.5458526573172258   0.7212285504135799   0.31836838938694273   0.5444391674984567   0.5263977915286694   0.12044953876186158   0.06874064240922237   0.6777197482290283   0.5127682853517493   0.5062675430152119   0.36271142353997643   0.3511762171667697   0.45336865926486336   0.1924460130141461   0.6973952819727792   0.9026019438374137   0.6166550453473159   0.4015291446153402   0.2854639532730119   0.4460744334521483   0.062232655525309793   0.5647408165750296   0.7407609764708422   0.44587164919581285   0.5163799982080841   0.8435122661614497   0.4223925870838994   0.9014324816973561   0.9899822066794147   0.7230627273995881   0.353651944674677   0.22371273346832787   0.4772139213276654   0.21679518438437617   0.9909405211347005   0.8725365163015582   0.02384526206280202   0.024349171370230068   0.2935452391619214   0.9699345724641445   0.4071902167154862   0.6228200267548898   0.008081285888909507   0.5238601390119961   0.3449575611901764   0.058079210179860154   0.2673203094180674   0.07798848981618331   0.8285775629820923   0.21456694401841042   0.844927722334168   0.17655600811882716   0.8385953563026777   0.49150421661882226   0.49127577765949104   0.9528432746504993   0.3613814349750123   0.2747090322344461   0.5003352565247905   0.08030675834894116   0.3375361729122103   0.250359860864216
0.20679001736286906   0.11037218588479669   0.9303459561967241   0.6275398341093262   0.19870873147395954   0.5865120468728006   0.5853883950065476   0.5694606239294661   0.9313884220558921   0.5085235570566172   0.7568108320244553   0.35489367991105564   0.08646069972172413   0.33196754893779007   0.9182154757217776   0.8633894632922333   0.5951849220622331   0.3791242742872908   0.5568340407467653   0.5886804310577872   0.09484966553744263   0.2988175159383496   0.21929786783455507   0.3383205701935712   0.8880596481745736   0.18844533005355293   0.288951911637831   0.710780736084245   0.689350916700614   0.6019332831807523   0.7035635166312834   0.14132011215477894   0.7579624946447219   0.09340972612413513   0.946752684606828   0.7864264322437233   0.6715017949229978   0.7614421771863451   0.028537208885050448   0.92303696895149   0.07631687286076466   0.38231790289905426   0.4717031681382851   0.33435653789370273   0.981467207323322   0.08350038696070466   0.25240530030373004   0.9960359677001315   0.09340755914874846   0.8950550569071517   0.963453388665899   0.28525523161588645   0.40405664244813444   0.29312177372639936   0.25988987203461567   0.1439351194611075   0.6460941478034126   0.19971204760226424   0.31313718742778757   0.3575086872173842   0.9745923528804148   0.4382698704159192   0.2845999785427371   0.43447171826589426
0.8982754800196502   0.05595196751686489   0.812896810404452   0.10011518037219154   0.9168082726963281   0.9724515805561602   0.560491510100722   0.10407921267206005   0.8234007135475797   0.07739652364900848   0.5970381214348229   0.8188239810561736   0.4193440710994452   0.7842747499226091   0.3371482494002073   0.6748888615950661   0.7732499232960327   0.5845627023203449   0.02401106197241974   0.31738017437768185   0.7986575704156178   0.1462928319044257   0.7394110834296826   0.8829084561117876   0.9003820903959677   0.09034086438756082   0.9265142730252306   0.7827932757395961   0.9835738176996396   0.1178892838314006   0.36602276292450864   0.678714063067536   0.16017310415205993   0.04049276018239211   0.7689846414896857   0.8598900820113624   0.7408290330526147   0.25621801025978297   0.4318363920894784   0.18500122041629638   0.967579109756582   0.6716553079394381   0.4078253301170586   0.8676210460386146   0.16892153934096418   0.5253624760350124   0.668414246687376   0.9847125899268269   0.2685394489449965   0.43502161164745157   0.7418999736621454   0.2019193141872308   0.2849656312453569   0.31713232781605094   0.3758772107376368   0.5232052511196947   0.12479252709329697   0.2766395676336589   0.6068925692479511   0.6633151691083323   0.38396349404068225   0.02042155737387586   0.17505617715847277   0.478313948692036
0.41638438428410024   0.34876624943443774   0.7672308470414142   0.6106929026534215   0.24746284494313603   0.8234037733994254   0.09881660035403815   0.6259803127265945   0.9789233959981395   0.3883821617519738   0.3569166266918927   0.42406099853936374   0.6939577647527826   0.07124983393592284   0.9810394159542559   0.9008557474196689   0.5691652376594857   0.794610266302264   0.3741468467063048   0.23754057831133663   0.1852017436188034   0.7741887089283881   0.19909066954783208   0.7592266296193007   0.7688173593347032   0.42542245949395036   0.4318598225064179   0.14853372696587924   0.5213545143915671   0.602018686094525   0.3330432221523798   0.5225534142392847   0.5424311183934276   0.21363652434255118   0.9761265954604871   0.098492415699921   0.848473353640645   0.14238669040662835   0.995087179506231   0.19763666828025206   0.27930811598115934   0.3477764241043644   0.6209403327999262   0.9600960899689155   0.09410637236235594   0.5735877151759762   0.42184966325209416   0.20086946034961478   0.3252890130276528   0.14816525568202588   0.9899898407456762   0.05233573338373553   0.8039344986360857   0.5461465695875009   0.6569466185932965   0.5297823191444508   0.261503380242658   0.33251004524494965   0.6808200231328094   0.43128990344452983   0.41303002660201305   0.19012335483832132   0.6857328436265784   0.23365323516427777
0.1337219106208537   0.842346930733957   0.06479251082665212   0.27355714519536234   0.03961553825849776   0.2687592155579807   0.642942847574558   0.07268768484574756   0.7143265252308449   0.12059395987595488   0.6529530068288817   0.02035195146201202   0.9103920265947594   0.574447390288454   0.9960063882355853   0.4905696323175612   0.6488886463521013   0.24193734504350434   0.3151863651027758   0.05927972887303137   0.23585861975008832   0.05181399020518301   0.6294535214761975   0.8256264937087536   0.10213670912923462   0.20946705947122604   0.5646610106495453   0.5520693485133913   0.06252117087073686   0.9407078439132452   0.9217181630749873   0.47938166366764373   0.3481946456398919   0.8201138840372905   0.26876515624610564   0.4590297122056317   0.4378026190451325   0.24566649374883642   0.2727587680105204   0.9684600798880705   0.7889139726930312   0.003729148705332078   0.9575724029077446   0.9091803510150391   0.5530553529429428   0.9519151585001491   0.32811888143154716   0.08355385730628553   0.4509186438137083   0.7424480990289231   0.7634578707820018   0.5314845087928942   0.3883974729429714   0.8017402551156777   0.8417397077070145   0.052102845125250555   0.04020282730307951   0.9816263710783873   0.5729745514609088   0.5930731329196188   0.6024002082579469   0.7359598773295509   0.3002157834503884   0.6246130530315483
0.8134862355649158   0.7322307286242188   0.3426433805426438   0.7154327020165092   0.26043088262197295   0.7803155701240697   0.014524499111096652   0.6318788447102237   0.8095122388082647   0.03786747109514672   0.2510666283290948   0.10039433591732945   0.4211147658652933   0.23612721597946898   0.40932692062208037   0.0482914907920789   0.3809119385622138   0.25450084490108166   0.8363523691611716   0.45521835787246007   0.7785117303042668   0.5185409675715308   0.5361365857107832   0.8306053048409117   0.965025494739351   0.786310238947312   0.19349320516813936   0.11517260282440243   0.7045946121173781   0.005994668823242197   0.1789687060570427   0.48329375811417874   0.8950823733091134   0.9681271977280955   0.9279020777279479   0.38289942219684925   0.4739676074438201   0.7319999817486265   0.5185751571058675   0.33460793140477035   0.09305566888160634   0.47749913684754486   0.6822227879446959   0.8793895735323103   0.31454393857733953   0.9589581692760141   0.14608620223391278   0.048784268691398645   0.3495184438379886   0.17264793032870213   0.9525929970657734   0.9336116658669962   0.6449238317206105   0.16665326150545992   0.7736242910087306   0.4503179077528175   0.7498414584114971   0.19852606377736443   0.8457222132807828   0.06741848555596823   0.27587385096767697   0.4665260820287379   0.3271470561749153   0.7328105541511979
0.18281818208607065   0.989026945181193   0.6449242682302193   0.8534209806188876   0.8682742435087311   0.03006877590517904   0.4988380659963066   0.8046367119274889   0.5187557996707426   0.8574208455764769   0.5462450689305332   0.8710250460604927   0.8738319679501321   0.690767584071017   0.7726207779218025   0.4207071383076752   0.12399050953863497   0.4922415202936526   0.9268985646410196   0.35328865275170696   0.848116658570958   0.025715438264914632   0.5997515084661044   0.6204780986005091   0.6652984764848874   0.03668849308372153   0.9548272402358849   0.7670571179816216   0.7970242329761562   0.006619717178542492   0.4559891742395784   0.9624204060541326   0.2782684333054137   0.14919887160206557   0.9097441053090453   0.09139535999363994   0.4044364653552816   0.45843128753104856   0.1371233273872428   0.6706882216859648   0.2804459558166466   0.966189767237396   0.21022476274622318   0.3173995689342578   0.43232929724568864   0.9404743289724814   0.6104732542801188   0.6969214703337487   0.7670308207608013   0.9037858358887598   0.6556460140442338   0.9298643523521272   0.9700065877846451   0.8971661187102173   0.1996568398046554   0.9674439462979946   0.6917381544792315   0.7479672471081518   0.2899127344956101   0.8760485863043547   0.2873016891239498   0.2895359595771032   0.1527894071083673   0.20536036461838988
0.006855733307303231   0.3233461923397072   0.9425646443621442   0.8879607956841321   0.5745264360616146   0.38287186336722584   0.3320913900820253   0.19103932535038334   0.8074956153008133   0.479086027478466   0.6764453760377914   0.26117497299825615   0.8374890275161682   0.5819199087682487   0.47678853623313605   0.2937310267002616   0.14575087303693676   0.833952661660097   0.18687580173752597   0.4176824403959069   0.858449183912987   0.5444167020829938   0.03408639462915865   0.21232207577751705   0.8515934506056837   0.22107050974328651   0.09152175026701452   0.324361280093385   0.27706701454406907   0.8381986463760607   0.7594303601849892   0.13332195474300165   0.4695713992432558   0.3591126188975946   0.08298498414719772   0.8721469817447455   0.6320823717270876   0.777192710129346   0.6061964479140617   0.578415955044484   0.48633149869015085   0.943240048469249   0.4193206461765357   0.16073351464857705   0.6278823147771639   0.39882334638625533   0.38523425154737706   0.94841143887106   0.7762888641714802   0.17775283664296881   0.2937125012803625   0.624050158777675   0.4992218496274111   0.33955419026690814   0.5342821410953733   0.4907282040346734   0.02965045038415533   0.9804415713693135   0.4512971569481756   0.6185812222899278   0.3975680786570677   0.20324886123996758   0.8451007090341139   0.040165267245443885
0.9112365799669169   0.2600088127707186   0.42578006285757825   0.8794317525968668   0.283354265189753   0.8611854663844632   0.0405458113102012   0.9310203137258068   0.5070654010182728   0.6834326297414944   0.7468333100298387   0.3069701549481318   0.007843551390861615   0.3438784394745863   0.21255116893446532   0.8162419509134584   0.9781931010067063   0.36343686810527276   0.7612540119862897   0.1976607286235306   0.5806250223496385   0.16018800686530515   0.9161533029521758   0.15749546137808673   0.6693884423827217   0.9001791940945866   0.49037324009459754   0.2780637087812199   0.3860341771929687   0.03899372771012335   0.44982742878439635   0.34704339505541304   0.8789687761746959   0.3555610979686289   0.7029941187545576   0.04007324010728123   0.8711252247838344   0.011682658494042653   0.49044294982009234   0.22383128919382278   0.892932123777128   0.64824579038877   0.7291889378338027   0.02617056057029218   0.31230710142748946   0.4880577835234648   0.8130356348816269   0.8686750991922054   0.6429186590447679   0.5878785894288782   0.3226623947870293   0.5906113904109855   0.25688448185179913   0.5488848617187548   0.872834966002633   0.24356799535557253   0.3779157056771032   0.19332376375012592   0.1698408472480753   0.2034947552482913   0.5067904808932688   0.18164110525608326   0.679397897427983   0.9796634660544685
0.6138583571161408   0.5333953148673133   0.9502089595941803   0.9534929054841763   0.3015512556886513   0.04533753134384857   0.13717332471255347   0.08481780629197087   0.6586325966438835   0.4574589419149704   0.8145109299255242   0.4942064158809853   0.4017481147920844   0.9085740801962155   0.9416759639228912   0.25063842052541274   0.023832409114981197   0.7152503164460896   0.7718351166748159   0.047143665277121466   0.5170419282217124   0.5336092111900064   0.09243721924683294   0.06748019922265294   0.9031835711055715   0.00021389632269306334   0.14222825965265262   0.1139872937384766   0.6016323154169202   0.9548763649788445   0.0050549349400991405   0.02916948744650572   0.9429997187730367   0.4974174230638741   0.19054400501457497   0.5349630715655204   0.5412516039809523   0.5888433428676585   0.24886804109168378   0.2843246510401077   0.5174191948659711   0.8735930264215689   0.4770329244168679   0.23718098576298619   0.0003772666442587349   0.33998381523156246   0.38459570517003494   0.16970078654033324   0.09719369553868723   0.33976991890886943   0.2423674455173823   0.05571349280185665   0.49556138012176704   0.3848935539300249   0.23731251057728317   0.026544005355350925   0.5525616613487304   0.8874761308661508   0.04676850556270819   0.49158093378983053   0.011310057367778136   0.2986327879984923   0.7979004644710244   0.20725628274972285
0.4938908625018071   0.4250397615769234   0.3208675400541565   0.9700752969867367   0.49351359585754834   0.08505594634536094   0.9362718348841216   0.8003745104464034   0.3963199003188611   0.7452860274364915   0.6939043893667394   0.7446610176445467   0.900758520197094   0.36039247350646664   0.4565918787894562   0.7181170122891959   0.34819685884836366   0.4729163426403158   0.409823373226748   0.22653607849936536   0.33688680148058553   0.17428355464182352   0.6119229087557235   0.01927979574964249   0.8429959389787784   0.7492437930649001   0.291055368701567   0.04920449876290582   0.3494823431212301   0.6641878467195391   0.3547835338174454   0.2488299883165024   0.9531624428023691   0.9189018192830476   0.6608791444507061   0.5041689706719557   0.052403922605274954   0.558509345776581   0.2042872656612499   0.7860519583827598   0.7042070637569113   0.08559300313626521   0.7944638924345019   0.5595158798833945   0.3673202622763258   0.9113094484944417   0.18254098367877838   0.5402360841337519   0.5243243232975473   0.16206565542954157   0.8914856149772113   0.4910315853708461   0.17484198017631722   0.4978778087100024   0.5367020811597659   0.24220159705434371   0.22167953737394822   0.5789759894269548   0.8758229367090599   0.7380326263823881   0.16927561476867325   0.020466643650373786   0.67153567104781   0.9519806679996283
0.465068551011762   0.9348736405141086   0.8770717786133081   0.39246478811623386   0.09774828873543617   0.02356419201966689   0.6945307949345297   0.852228703982482   0.5734239654378889   0.8614985365901253   0.8030451799573183   0.36119711861163584   0.3985819852615716   0.3636207278801229   0.26634309879755236   0.11899552155729212   0.17690244788762338   0.7846447384531681   0.3905201620884925   0.38096289517490406   0.007626833118950135   0.7641780948027943   0.7189844910406825   0.42898222717527573   0.5425582821071882   0.8293044542886857   0.8419127124273744   0.036517439059041826   0.44480999337175203   0.8057402622690188   0.14738191749284474   0.18428873507655988   0.8713860279338632   0.9442417256788935   0.3443367375355264   0.823091616464924   0.47280404267229154   0.5806209977987706   0.07799363873797403   0.7040960949076319   0.29590159478466815   0.7959762593456026   0.6874734766494816   0.32313319973272786   0.288274761665718   0.03179816454280826   0.968488985608799   0.8941509725574521   0.7457164795585298   0.20249371025412252   0.12657627318142467   0.8576335334984103   0.30090648618677784   0.3967534479851037   0.9791943556885799   0.6733447984218505   0.4295204582529147   0.4525117223062102   0.6348576181530535   0.8502531819569265   0.9567164155806231   0.8718907245074395   0.5568639794150795   0.1461570870492945
0.660814820795955   0.07591446516183695   0.8693905027655979   0.8230238873165666   0.3725400591302369   0.044116300619028694   0.9009015171567989   0.9288729147591145   0.6268235795717071   0.8416225903649062   0.7743252439753742   0.07123938126070412   0.3259170933849292   0.44486914237980246   0.7951308882867942   0.39789458283885365   0.8963966351320145   0.9923574200735923   0.16027327013374074   0.5476414008819273   0.9396802195513915   0.12046669556615279   0.6034092907186612   0.4014843138326327   0.2788653987554365   0.04455223040431584   0.7340187879530633   0.5784604265160661   0.9063253396251996   0.0004359297852871483   0.8331172707962645   0.6495875117569516   0.2795017600534925   0.15881333942038098   0.0587920268208903   0.5783481304962474   0.9535846666685632   0.7139441970405785   0.26366113853409606   0.18045354765739385   0.05718803153654874   0.7215867769669863   0.10338786840035531   0.6328121467754666   0.11750781198515732   0.6011200814008334   0.49997857768169407   0.23132783294283393   0.8386424132297209   0.5565678509965176   0.7659597897286308   0.6528674064267679   0.9323170736045213   0.5561319212112305   0.9328425189323662   0.0032798946698162374   0.6528153135510287   0.39731858179084945   0.874050492111476   0.42493176417356876   0.6992306468824655   0.6833743847502709   0.6103893535773799   0.24447821651617488
0.6420426153459168   0.9617876077832848   0.5070014851770246   0.6116660697407083   0.5245348033607594   0.3606675263824513   0.007022907495330553   0.3803382367978743   0.6858923901310386   0.8040996753859337   0.2410631177666998   0.7274708303711065   0.7535753165265173   0.2479677541747033   0.30822059883433356   0.7241909357012902   0.10076000297548852   0.8506491723838538   0.43417010672285755   0.2992591715277215   0.40152935609302304   0.16727478763358292   0.8237807531454776   0.05478095501154661   0.7594867407471063   0.2054871798502982   0.316779267968453   0.44311488527083837   0.23495193738634684   0.8448196534678469   0.30975636047312244   0.06277664847296402   0.5490595472553083   0.0407199780819132   0.06869324270642264   0.33530581810185756   0.7954842307287909   0.7927522239072099   0.7604726438720891   0.6111148824005673   0.6947242277533024   0.942103051523356   0.3263025371492316   0.3118557108728458   0.2931948716602794   0.7748282638897731   0.5025217840037539   0.2570747558612992   0.5337081309131732   0.5693410840394749   0.18574251603530093   0.8139598705904608   0.2987561935268263   0.724521430571628   0.8759861555621785   0.7511832221174968   0.749696646271518   0.6838014524897148   0.8072929128557558   0.4158774040156393   0.9542124155427271   0.8910492285825049   0.046820268983666716   0.804762521615072
0.2594881877894247   0.9489461770591489   0.7205177318344351   0.4929068107422262   0.9662933161291453   0.1741179131693757   0.2179959478306812   0.235832054880927   0.43258518521597217   0.6047768291299008   0.032253431795380295   0.4218721842904662   0.13382899168914586   0.8802553985582727   0.1562672762332018   0.6706889621729694   0.3841323454176278   0.19645394606855798   0.348974363377446   0.2548115581573301   0.42991992987490074   0.3054047174860531   0.30215409439377927   0.45004903654225814   0.17043174208547607   0.3564585404269043   0.5816363625593441   0.9571422258000319   0.2041384259563308   0.18234062725752856   0.3636404147286629   0.7213101709191049   0.7715532407403587   0.5775637981276278   0.3313869829332826   0.29943798662863874   0.6377242490512128   0.697308399569355   0.17511970670008078   0.6287490244556694   0.25359190363358497   0.500854453500797   0.8261453433226348   0.37393746629833924   0.8236719737586843   0.19544973601474394   0.5239912489288555   0.9238884297560811   0.6532402316732082   0.8389911955878396   0.9423548863695114   0.9667462039560492   0.44910180571687736   0.6566505683303111   0.5787144716408485   0.24543603303694422   0.6775485649765187   0.07908677020268332   0.2473274887075659   0.9459980464083055   0.039824315925305886   0.3817783706333283   0.07220778200748512   0.31724902195263616
0.7862324122917209   0.8809239171325313   0.2460624386848503   0.9433115556542969   0.9625604385330366   0.6854741811177874   0.7220711897559948   0.01942312589821582   0.30932020685982853   0.8464829855299476   0.7797163033864833   0.05267692194216666   0.8602184011429511   0.1898324171996365   0.20100183174563485   0.8072408889052224   0.18266983616643245   0.11074564699695318   0.953674343038069   0.861242842496917   0.14284552024112657   0.7289672763636249   0.8814665610305839   0.5439938205442808   0.35661310794940565   0.8480433592310936   0.6354041223457335   0.6006822648899839   0.39405266941636896   0.16256917811330635   0.9133329325897387   0.5812591389917681   0.08473246255654047   0.31608619258335874   0.13361662920325537   0.5285822170496014   0.22451406141358932   0.12625377538372223   0.9326147974576205   0.7213413281443789   0.04184422524715688   0.015508128386769052   0.9789404544195516   0.860098485647462   0.8989987050060303   0.28654085202314417   0.09747389338896773   0.31610466510318125   0.5423855970566247   0.4384974927920505   0.4620697710432342   0.7154224002131974   0.14833292764025569   0.2759283146787442   0.5487368384534955   0.13416326122142938   0.06360046508371521   0.9598421220953854   0.4151202092502401   0.605581044171828   0.8390864036701259   0.8335883467116633   0.4825054117926196   0.8842397160274491
0.797242178422969   0.8180802183248942   0.5035649573730681   0.024141230379987045   0.8982434734169387   0.53153936630175   0.4060910639841003   0.7080365652768058   0.355857876360314   0.09304187350969947   0.9440212929408661   0.9926141650636083   0.20752494872005833   0.8171135588309553   0.3952844544873706   0.858450903842179   0.14392448363634314   0.8572714367355698   0.9801642452371305   0.252869859670351   0.30483807996621726   0.023683090023906634   0.4976588334445109   0.3686301436429019   0.5075959015432483   0.20560287169901248   0.9940938760714428   0.3444889132629149   0.6093524281263095   0.6740635053972625   0.5880028120873426   0.6364523479861091   0.25349455176599556   0.581021631887563   0.6439815191464765   0.6438381829225007   0.04596960304593722   0.7639080730566077   0.2486970646591059   0.7853872790803217   0.9020451194095941   0.9066366363210379   0.2685328194219754   0.5325174194099707   0.5972070394433768   0.8829535462971312   0.7708739859774645   0.16388727576706877   0.08961113790012858   0.6773506745981187   0.7767801099060215   0.8193983625041539   0.480258709773819   0.003287169200856278   0.188777297818679   0.18294601451804476   0.22676415800782346   0.42226553731329325   0.5447957786722025   0.5391078315955441   0.18079455496188623   0.6583574642566855   0.29609871401309656   0.7537205525152224
0.27874943555229215   0.7517208279356477   0.027565894591121184   0.22120313310525166   0.6815423961089153   0.8687672816385165   0.2566919086136567   0.0573158573381829   0.5919312582087868   0.19141660704039773   0.4799117987076351   0.23791749483402905   0.11167254843496774   0.18812943783954145   0.29113450088895615   0.05497148031598427   0.8849083904271443   0.7658639005262482   0.7463387222167537   0.5158636487204402   0.7041138354652581   0.1075064362695626   0.45024000820365706   0.7621430962052179   0.4253643999129659   0.35578560833391487   0.4226741136125359   0.5409399630999662   0.7438220038040506   0.4870183266953984   0.1659822049988792   0.48362410576178333   0.1518907455952638   0.2956017196550007   0.686070406291244   0.24570661092775425   0.04021819716029607   0.10747228181545927   0.39493590540228796   0.19073513061177   0.15530980673315178   0.3416083812892111   0.6485971831855343   0.6748714818913297   0.45119597126789374   0.2341019450196485   0.1983571749818772   0.9127283856861119   0.02583157135492785   0.8783163366857336   0.7756830613693413   0.3717884225861457   0.2820095675508773   0.3912980099903352   0.6097008563704621   0.8881643168243624   0.13011882195561347   0.09569629033533447   0.9236304500792181   0.6424577058966081   0.0899006247953174   0.9882240085198752   0.5286945446769301   0.4517225752848381
0.9345908180621656   0.6466156272306641   0.8800973614913958   0.7768510933935083   0.48339484679427186   0.4125136822110156   0.6817401865095186   0.8641227077073964   0.457563275439344   0.534197345525282   0.9060571251401773   0.49233428512125077   0.17555370788846672   0.1428993355349468   0.2963562687697152   0.6041699682968884   0.04543488593285327   0.04720304519961234   0.37272581869049715   0.9617122624002802   0.9555342611375359   0.05897903667973713   0.844031274013567   0.5099896871154421   0.020943443075370275   0.412363409449073   0.9639339125221712   0.7331385937219337   0.5375485962810984   0.9998497272380574   0.2821937260126525   0.8690158860145373   0.0799853208417544   0.46565238171277545   0.3761366008724752   0.3766816008932865   0.9044316129532877   0.32275304617782863   0.07978033210275995   0.7725116325963981   0.8589967270204344   0.2755500009782163   0.7070545134122628   0.8107993701961179   0.9034624658828985   0.21657096429847916   0.8630232393986957   0.30080968308067585   0.8825190228075283   0.8042075548494061   0.8990893268765245   0.5676710893587421   0.34497042652642984   0.8043578276113487   0.6168956008638721   0.6986552033442048   0.2649851056846754   0.33870544589857327   0.24075899999139688   0.3219736024509184   0.36055349273138776   0.01595239972074461   0.16097866788863693   0.5494619698545202
0.5015567657109534   0.7404023987425283   0.45392415447637413   0.7386625996584023   0.5980942998280548   0.5238314344440491   0.5909009150776784   0.4378529165777264   0.7155752770205266   0.719623879594643   0.6918115882011538   0.8701818272189843   0.3706048504940968   0.9152660519832942   0.07491598733728176   0.1715266238747794   0.10561974480942136   0.576560606084721   0.8341569873458848   0.849553021423861   0.7450662520780336   0.5606082063639765   0.6731783194572479   0.30009105156934085   0.24350948636708022   0.8202058076214481   0.2192541649808738   0.5614284519109386   0.6454151865390253   0.296374373177399   0.6283532499031954   0.12357553533321215   0.9298399095184987   0.576750493582756   0.9365416617020416   0.25339370811422784   0.559235059024402   0.6614844415994617   0.8616256743647598   0.08186708423944845   0.4536153142149805   0.08492383551474067   0.027468687018874942   0.2323140628155874   0.7085490621369469   0.5243156291507642   0.35429036756162696   0.9322230112462465   0.46503957576986676   0.7041098215293161   0.13503620258075316   0.37079455933530797   0.8196243892308414   0.4077354483519171   0.5066829526775578   0.24721902400209583   0.8897844797123426   0.8309849547691611   0.5701412909755161   0.9938253158878679   0.3305494206879408   0.16950051316969938   0.7085156166107563   0.9119582316484195
0.8769341064729602   0.08457667765495872   0.6810469295918814   0.6796441688328321   0.16838504433601326   0.5602610485041944   0.3267565620302544   0.7474211575865856   0.7033454685661465   0.8561512269748784   0.19172035944950122   0.3766265982512776   0.8837210793353051   0.4484157786229613   0.6850374067719435   0.12940757424918173   0.9939365996229624   0.6174308238538002   0.11489611579642732   0.13558225836131377   0.6633871789350216   0.44793031068410083   0.406380499185671   0.22362402671289427   0.7864530724620614   0.36335363302914214   0.7253335695937896   0.5439798578800622   0.6180680281260482   0.8030925845249476   0.3985770075635352   0.7965587002934766   0.9147225595599017   0.9469413575500693   0.20685664811403398   0.41993210204219905   0.031001480224596558   0.4985255789271079   0.5218192413420905   0.29052452779301735   0.03706488060163414   0.8810947550733077   0.4069231255456632   0.15494226943170356   0.3736777016666125   0.4331644443892069   0.000542626359992191   0.9313182427188093   0.5872246292045511   0.06981081136006478   0.2752090567662026   0.3873383848387471   0.9691566010785029   0.26671822683511714   0.8766320492026674   0.5907796845452705   0.05443404151860125   0.3197768692850479   0.6697754010886334   0.17084758250307142   0.02343256129400469   0.82125129035794   0.1479561597465429   0.8803230547100541
0.9863676806923706   0.9401565352846323   0.7410330342008797   0.7253807852783505   0.6126899790257581   0.5069920908954253   0.7404904078408875   0.7940625425595412   0.025465349821206972   0.43718127953536057   0.46528135107468493   0.4067241577207941   0.05630874874270407   0.1704630527002434   0.5886493018720176   0.8159444731755237   0.0018747072241028216   0.8506861834151955   0.9188739007833842   0.6450968906724522   0.9784421459300982   0.02943489305725551   0.7709177410368413   0.7647738359623982   0.9920744652377276   0.08927835777262327   0.02988470683596155   0.03939305068404768   0.3793844862119695   0.582286266877198   0.289394298995074   0.24533050812450644   0.35391913639076256   0.14510498734183738   0.8241129479203891   0.8386063504037123   0.29761038764805847   0.974641934641594   0.23546364604837153   0.02266187722818862   0.29573568042395565   0.12395575122639849   0.31658974526498734   0.37756498655573634   0.31729353449385755   0.09452085816914298   0.5456720042281461   0.6127911505933381   0.32521906925613   0.005242500396519708   0.5157872973921845   0.5733980999092905   0.9458345830441605   0.42295623351932177   0.22639299839711052   0.328067591784784   0.5919154466533979   0.2778512461774844   0.40228005047672144   0.4894612413810717   0.2943050590053394   0.3032093115358904   0.1668164044283499   0.4667993641528831
0.9985693785813837   0.17925356030949197   0.8502266591633626   0.08923437759714677   0.6812758440875262   0.08473270214034898   0.30455465493521644   0.4764432270038086   0.3560567748313962   0.07949020174382927   0.788767357543032   0.9030451270945181   0.41022219178723573   0.6565339682245075   0.5623743591459214   0.5749775353097341   0.8183067451338379   0.3786827220470231   0.16009430866919996   0.08551629392866238   0.5240016861284985   0.07547341051113264   0.99327790424085   0.6187169297757793   0.5254323075471149   0.8962198502016406   0.14305124507748748   0.5294825521786325   0.8441564634595887   0.8114871480612917   0.8384965901422711   0.05303932517482388   0.4880996886281926   0.7319969463174625   0.04972923259923912   0.14999419808030573   0.07787749684095681   0.07546297809295495   0.48735487345331774   0.5750166627705716   0.2595707517071189   0.6967802560459319   0.3272605647841178   0.4895003688419093   0.7355690655786203   0.6213068455347992   0.33398266054326775   0.87078343906613   0.21013675803150547   0.7250869953331586   0.19093141546578024   0.3413008868874975   0.3659802945719167   0.9135998472718668   0.3524348253235092   0.28826156171267364   0.8778806059437242   0.18160290095440443   0.3027055927242701   0.13826736363236788   0.8000031091027674   0.10613992286144946   0.8153507192709524   0.5632507008617963
0.5404323573956484   0.4093596668155176   0.48809015448683457   0.07375033201988698   0.8048632918170281   0.7880528212807184   0.15410749394356685   0.20296689295375697   0.5947265337855226   0.06296582594755983   0.9631760784777866   0.8616660060662594   0.2287462392136059   0.14936597867569298   0.6107412531542774   0.5734044443535858   0.35086563326988174   0.9677630777212886   0.3080356604300073   0.435137080721218   0.5508625241671143   0.8616231548598391   0.4926849411590549   0.8718863798594217   0.01043016677146593   0.4522634880443215   0.004594786672220347   0.7981360478395347   0.20556687495443784   0.6642106667636031   0.8504872927286535   0.5951691548857777   0.6108403411689152   0.6012448408160433   0.8873112142508669   0.7335031488195183   0.38209410195530935   0.45187886214035033   0.27656996109658954   0.1600987044659324   0.031228468685427595   0.4841157844190618   0.9685343006665822   0.7249616237447145   0.4803659445183132   0.6224926295592227   0.4758493595075273   0.8530752438852928   0.4699357777468473   0.1702291415149012   0.471254572835307   0.054939196045758025   0.26436890279240943   0.5060184747512981   0.6207672801066535   0.45977004115998027   0.6535285616234943   0.9047736339352548   0.7334560658557866   0.726266892340462   0.2714344596681849   0.4528947717949045   0.45688610475919705   0.5661681878745296
0.24020599098275733   0.9687789873758427   0.4883518040926148   0.8412065641298151   0.7598400464644441   0.34628635781662004   0.0125024445850875   0.9881313202445223   0.28990426871759684   0.17605721630171883   0.5412478717497805   0.9331921241987643   0.025535365925187358   0.6700387415504208   0.9204805916431271   0.4734220830387841   0.37200680430169314   0.765265107615166   0.18702452578734055   0.747155190698322   0.1005723446335082   0.31237033582026147   0.7301384210281435   0.1809870028237925   0.8603663536507509   0.34359134844441874   0.24178661693552872   0.33978043869397734   0.10052630718630677   0.9973049906277988   0.2292841723504412   0.351649118449455   0.81062203846871   0.8212477743260799   0.6880363006006607   0.41845699425069066   0.7850866725435226   0.15120903277565914   0.7675557089575336   0.9450349112119065   0.41307986824182946   0.3859439251604932   0.580531183170193   0.19787972051358452   0.3125075236083213   0.07357358934023175   0.8503927621420495   0.016892717689792044   0.4521411699575704   0.729982240895813   0.6086061452065208   0.6771122789958147   0.35161486277126364   0.7326772502680143   0.37932197285607955   0.3254631605463597   0.5409928243025537   0.9114294759419344   0.6912856722554189   0.9070061662956691   0.7559061517590311   0.7602204431662752   0.9237299632978853   0.9619712550837625
0.34282628351720157   0.37427651800578204   0.3431987801276923   0.764091534570178   0.030318759908880295   0.30070292866555026   0.4928060179856428   0.7471988168803859   0.5781775899513099   0.5707206877697373   0.884199872779122   0.07008653788457123   0.22656272718004625   0.8380434375017229   0.5048778999230424   0.7446233773382115   0.6855699028774925   0.9266139615597886   0.8135922276676236   0.8376172110425425   0.9296637511184614   0.16639351839351332   0.8898622643697383   0.8756459559587799   0.5868374676012599   0.7921170003877313   0.546663484242046   0.11155442138860201   0.5565187076923797   0.491414071722181   0.05385746625640324   0.3643556045082161   0.9783411177410697   0.9206933839524437   0.16965759347728124   0.2942690666236449   0.7517783905610235   0.08264994645072073   0.6647796935542387   0.5496456892854333   0.06620848768353092   0.15603598489093215   0.8511874658866152   0.7120284782428908   0.13654473656506944   0.9896424664974188   0.9613252015168768   0.8363825222841109   0.5497072689638095   0.19752546610968758   0.41466171727483087   0.7248281008955089   0.9931885612714298   0.7061113943875066   0.3608042510184276   0.3604724963872928   0.014847443530360155   0.7854180104350629   0.19114665754114638   0.06620342976364794   0.26306905296933664   0.7027680639843421   0.5263669639869076   0.5165577404782146
0.19686056528580573   0.54673207909341   0.6751794981002924   0.8045292622353237   0.06031582872073631   0.5570896125959911   0.7138542965834156   0.9681467399512128   0.5106085597569268   0.3595641464863036   0.29919257930858467   0.24331863905570394   0.5174199984854969   0.6534527520987969   0.9383883282901571   0.8828461426684111   0.5025725549551368   0.8680347416637341   0.7472416707490107   0.8166427129047632   0.2395035019858001   0.16526667767939193   0.22087470676210308   0.3000849724265486   0.042642936699994353   0.6185345985859819   0.5456952086618106   0.49555571019122485   0.982327107979258   0.061444985989990805   0.8318409120783951   0.527408970240012   0.4717185482223312   0.7018808395036873   0.5326483327698104   0.2840903311843081   0.9542985497368344   0.048428087404890276   0.5942600044796533   0.401244188515897   0.45172599478169756   0.18039334574115617   0.8470183337306426   0.5846014756111337   0.21222249279589747   0.01512666806176425   0.6261436269685395   0.2845165031845852   0.1695795560959031   0.3965920694757823   0.08044841830672891   0.7889607929933603   0.18725244811664507   0.3351470834857915   0.24860750622833383   0.2615518227533483   0.7155338998943138   0.6332662439821043   0.7159591734585234   0.9774614915690402   0.7612353501574796   0.5848381565772139   0.12169916897887015   0.5762173030531432
0.30950935537578195   0.40444481083605777   0.2746808352482275   0.9916158274420095   0.09728686257988449   0.38931814277429355   0.648537208279688   0.7070993242574243   0.9277073064839814   0.9927260732985113   0.5680887899729591   0.918138531264064   0.7404548583673363   0.6575789898127198   0.3194812837446252   0.6565867085107157   0.024920958473022437   0.024312745830615497   0.6035221102861017   0.6791252169416754   0.2636856083155429   0.43947458925340155   0.48182294130723163   0.1029079138885322   0.9541762529397609   0.03502977841734374   0.2071421060590041   0.11129208644652275   0.8568893903598764   0.6457116356430502   0.5586048977793161   0.4041927621890985   0.9291820838758951   0.652985562344539   0.9905161078063571   0.4860542309250346   0.18872722550855878   0.9954065725318192   0.6710348240617319   0.829467522414319   0.16380626703553636   0.9710938267012037   0.06751271377563012   0.15034230547264354   0.9001206587199935   0.5316192374478023   0.5856897724683985   0.047434391584111335   0.9459444057802325   0.4965894590304585   0.3785476664093944   0.9361423051375886   0.08905501542035606   0.8508778233874082   0.8199427686300783   0.5319495429484901   0.15987293154446097   0.19789226104286928   0.8294266608237212   0.0458953120234555   0.9711457060359022   0.20248568851105006   0.15839183676198934   0.21642778960913653
0.8073394390003659   0.2313918618098463   0.09087912298635922   0.06608548413649301   0.9072187802803724   0.6997726243620441   0.5051893505179608   0.01865109255238167   0.9612743745001399   0.20318316533158565   0.1266416841085663   0.08250878741479309   0.8722193590797839   0.35230534194417734   0.306698915478488   0.550559244466303   0.7123464275353228   0.1544130809013081   0.4772722546547668   0.5046639324428475   0.7412007214994206   0.951927392390258   0.31888041789277743   0.28823614283371096   0.9338612824990548   0.7205355305804118   0.2280012949064182   0.22215065869721795   0.02664250221868241   0.020762906218367596   0.7228119443884575   0.2034995661448363   0.06536812771854252   0.817579740886782   0.5961702602798912   0.1209907787300432   0.19314876863875868   0.4652743989426046   0.2894713448014032   0.5704315342637402   0.48080234110343584   0.3108613180412965   0.8121990901466364   0.0657676018208927   0.7396016196040152   0.3589339256510385   0.493318672253859   0.7775314589871817   0.8057403371049604   0.6383983950706268   0.26531737734744076   0.5553808002899637   0.7790978348862779   0.6176354888522592   0.5425054329589832   0.3518812341451275   0.7137297071677354   0.8000557479654772   0.9463351726790921   0.23089045541508427   0.5205809385289768   0.33478134902287265   0.6568638278776888   0.6604589211513441
0.03977859742554092   0.023920030981576117   0.8446647377310524   0.5946913193304514   0.30017697782152575   0.6649861053305376   0.35134606547719344   0.8171598603432696   0.4944366407165654   0.026587710259910833   0.08602868812975266   0.26177906005330587   0.7153388058302874   0.40895222140765164   0.5435232551707694   0.9098978259081784   0.00160909866255198   0.6088964734421745   0.5971880824916773   0.6790073704930941   0.48102816013357524   0.2741151244193018   0.9403242546139885   0.01854844934175003   0.4412495627080343   0.25019509343772567   0.09565951688293609   0.42385713001129866   0.14107258488650856   0.585208988107188   0.7443134514057427   0.606697269668029   0.6466359441699432   0.5586212778472772   0.65828476327599   0.34491820961472314   0.9312971383396558   0.14966905643962555   0.11476150810522061   0.4350203837065447   0.9296880396771038   0.5407725829974511   0.5175734256135432   0.7560130132134506   0.44865987954352854   0.2666574585781494   0.5772491709995548   0.7374645638717006   0.007410316835494252   0.016462365140423714   0.4815896541166187   0.31360743386040196   0.8663377319489857   0.4312533770332357   0.737276202710876   0.706910164192373   0.21970178777904253   0.8726320991859585   0.07899143943488601   0.3619919545776498   0.28840464943938676   0.7229630427463329   0.9642299313296654   0.926971570871105
0.358716609762283   0.18219045974888176   0.44665650571612214   0.17095855765765447   0.9100567302187544   0.9155330011707324   0.8694073347165674   0.4334939937859539   0.9026464133832602   0.8990706360303087   0.3878176805999487   0.11988655992555192   0.03630868143427449   0.467817258997073   0.6505414778890727   0.41297639573317896   0.816606893655232   0.5951851598111145   0.5715500384541867   0.05098444115552913   0.5282022442158452   0.8722221170647816   0.6073201071245213   0.12401287028442404   0.1694856344535622   0.6900316573158999   0.16066360140839916   0.9530543126267695   0.25942890423480774   0.7744986561451674   0.2912562666918318   0.5195603188408157   0.35678249085154756   0.8754280201148588   0.9034385860918831   0.3996737589152638   0.3204738094172731   0.4076107611177857   0.25289710820281036   0.9866973631820848   0.5038669157620411   0.8124256013066712   0.6813470697486237   0.9357129220265558   0.975664671546196   0.9402034842418896   0.07402696262410237   0.8117000517421317   0.8061790370926337   0.25017182692598977   0.9133633612157032   0.8586457391153621   0.5467501328578259   0.47567317078082233   0.6221070945238715   0.3390854202745464   0.18996764200627836   0.6002451506659636   0.7186685084319884   0.9394116613592826   0.8694938325890053   0.19263438954817785   0.465771400229178   0.9527142981771978
0.36562691682696413   0.38020878824150667   0.7844243304805544   0.017001376150642046   0.3899622452807682   0.44000530399961707   0.710397367856452   0.20530132440851037   0.5837832081881345   0.18983347707362727   0.7970340066407487   0.34665558529314827   0.03703307533030854   0.7141603062928049   0.17492691211687733   0.007570165018601867   0.8470654333240302   0.11391515562684132   0.45625840368488896   0.06815850365931926   0.9775716007350249   0.9212807660786635   0.990487003455711   0.1154442054821215   0.6119446839080608   0.5410719778371568   0.2060626729751566   0.09844282933147946   0.22198243862729253   0.10106667383753976   0.4956653051187046   0.8931415049229691   0.638199230439158   0.9112331967639125   0.6986312984779558   0.5464859196298208   0.6011661551088495   0.19707289047110757   0.5237043863610785   0.538915754611219   0.7541007217848194   0.08315773484426625   0.06744598267618954   0.4707572509518997   0.7765291210497944   0.16187696876560279   0.07695897922047859   0.3553130454697782   0.16458443714173365   0.620804990928446   0.870896306245322   0.25687021613829875   0.9426019985144412   0.5197383170909062   0.3752310011266174   0.3637287112153296   0.3044027680752831   0.6085051203269938   0.6765997026486615   0.8172427915855088   0.7032366129664336   0.4114322298558862   0.1528953162875831   0.27832703697428984
0.9491358911816142   0.3282744950116199   0.08544933361139356   0.8075697860223902   0.17260677013181983   0.1663975262460171   0.008490354390914966   0.45225674055261195   0.008022332990086176   0.5455925353175711   0.13759404814559295   0.1953865244143132   0.06542033447564505   0.025854218226664904   0.7623630470189755   0.8316578131989836   0.761017566400362   0.4173490978996712   0.08576334437031395   0.01441502161347479   0.057780953433928396   0.005916868043785016   0.9328680280827308   0.736087984639185   0.10864506225231413   0.6776423730321651   0.8474186944713373   0.9285181986167949   0.9360382921204943   0.511244846786148   0.8389283400804223   0.4762614580641829   0.9280159591304081   0.9656523114685769   0.7013342919348293   0.2808749336498697   0.862595624654763   0.939798093241912   0.9389712449158538   0.4492171204508861   0.1015780582544011   0.5224489953422408   0.8532079005455399   0.4348020988374113   0.0437971048204727   0.5165321272984558   0.920339872462809   0.6987141141982264   0.9351520425681585   0.8388897542662906   0.07292117799147173   0.7701959155814315   0.9991137504476643   0.3276449074801427   0.2339928379110494   0.2939344575172486   0.07109779131725615   0.3619925960115658   0.53265854597622   0.013059523867378933   0.20850216666249308   0.4221945027696538   0.5936873010603662   0.5638424034164928
0.10692410840809198   0.8997455074274131   0.7404794005148263   0.12904030457908153   0.06312700358761929   0.3832133801289573   0.8201395280520173   0.4303261903808552   0.1279749610194607   0.5443236258626666   0.7472183500605456   0.6601302747994237   0.12886121057179645   0.21667871838252395   0.5132255121494962   0.3661958172821751   0.057763419254540295   0.8546861223709582   0.9805669661732761   0.35313629341479613   0.8492612525920472   0.43249161960130433   0.38687966511290994   0.7892938899983033   0.7423371441839552   0.5327461121738912   0.6464002645980836   0.6602535854192217   0.679210140596336   0.14953273204493397   0.8262607365460664   0.22992739503836657   0.5512351795768752   0.6052091061822673   0.07904238648552077   0.5697971202389429   0.4223739690050788   0.3885303877997434   0.5658168743360246   0.20360130295676782   0.36461054975053847   0.5338442654287853   0.5852499081627485   0.8504650095419717   0.5153492971584913   0.10135264582748095   0.19837024304983852   0.06117111954366838   0.7730121529745361   0.5686065336535897   0.5519699784517549   0.4009175341244466   0.09380201237820009   0.4190738016086557   0.7257092419056885   0.17099013908608002   0.5425668328013249   0.8138646954263884   0.6466668554201678   0.6011930188471372   0.12019286379624608   0.4253343076266449   0.08084998108414317   0.3975917158903693
0.7555823140457076   0.8914900421978597   0.4956000729213947   0.5471267063483977   0.24023301688721632   0.7901373963703787   0.2972298298715562   0.4859555868047293   0.4672208639126803   0.22153086271678907   0.7452598514198013   0.08503805268028264   0.37341885153448023   0.8024570611081333   0.019550609514112777   0.9140479135942026   0.8308520187331554   0.988592365681745   0.37288375409394503   0.31285489474706546   0.7106591549369092   0.5632580580551   0.2920337730098018   0.9152631788566962   0.9550768408912017   0.6717680158572403   0.7964337000884072   0.36813647250829856   0.7148438240039854   0.8816306194868616   0.499203870216851   0.8821808857035693   0.24762296009130505   0.6600997567700725   0.7539440187970496   0.7971428330232866   0.8742041085568248   0.8576426956619392   0.7343934092829368   0.883094919429084   0.04335208982366949   0.8690503299801943   0.36150965518899186   0.5702400246820185   0.3326929348867602   0.3057922719250942   0.06947588217919001   0.6549768458253223   0.37761609399555857   0.6340242560678538   0.27304218209078285   0.28684037331702383   0.6627722699915732   0.7523936365809922   0.7738383118739319   0.40465948761345455   0.41514930990026816   0.0922938798109197   0.019894293076882272   0.6075166545901679   0.5409452013434434   0.2346511841489805   0.2855008837939454   0.7244217351610839
0.49759311151977387   0.3656008541687863   0.9239912286049535   0.15418171047906534   0.16490017663301362   0.0598085822436921   0.8545153464257635   0.499204864653743   0.7872840826374551   0.4257843261758383   0.5814731643349806   0.2123644913367191   0.12451181264588185   0.673390689594846   0.8076348524610488   0.8077050037232646   0.7093625027456136   0.5810968097839263   0.7877405593841665   0.20018834913309666   0.16841730140217034   0.34644562563494585   0.5022396755902211   0.47576661397201275   0.6708241898823964   0.9808447714661596   0.5782484469852676   0.32158490349294744   0.5059240132493829   0.9210361892224674   0.723733100559504   0.8223800388392044   0.7186399306119278   0.4952518630466292   0.1422599362245233   0.6100155475024853   0.5941281179660459   0.8218611734517831   0.33462508376347455   0.8023105437792207   0.8847656152204323   0.24076436366785683   0.546884524379308   0.6021221946461242   0.7163483138182619   0.894318738032911   0.044644848789086936   0.12635558067411135   0.04552412393586545   0.9134739665667515   0.4663964018038194   0.8047706771811639   0.5396001106864826   0.992437777344284   0.7426633012443155   0.9823906383419595   0.8209601800745547   0.4971859142976548   0.6004033650197921   0.3723750908394741   0.22683206210850876   0.6753247408458717   0.2657782812563176   0.5700645470602533
0.34206644688807647   0.4345603771780148   0.7188937568770095   0.9679423524141293   0.6257181330698145   0.5402416391451038   0.6742489080879226   0.841586771740018   0.580194009133949   0.6267676725783523   0.2078525062841032   0.036816094558853964   0.04059389844746651   0.6343298952340684   0.4651892050397878   0.05442545621689449   0.21963371837291176   0.13714398093641353   0.8647858400199957   0.6820503653774204   0.992801656264403   0.46181924009054187   0.5990075587636781   0.11198581831716699   0.6507352093763266   0.027258862912527052   0.8801138018866685   0.14404346590303774   0.02501707630651201   0.48701722376742324   0.20586489379874598   0.30245669416301985   0.4448230671725629   0.8602495511890709   0.9980123875146427   0.26564059960416586   0.4042291687250964   0.22591965595500257   0.5328231824748549   0.21121514338727138   0.18459545035218466   0.08877567501858905   0.6680373424548592   0.5291647780098511   0.19179379408778166   0.6269564349280472   0.06902978369118118   0.41717895969268404   0.5410585847114551   0.5996975720155201   0.1889159818045126   0.2731354937896463   0.5160415084049431   0.11268034824809688   0.9830510880057667   0.9706787996266265   0.07121844123238018   0.252430797059026   0.9850387004911239   0.7050382000224605   0.6669892725072838   0.026511141104023413   0.4522155180162689   0.49382305663518916
0.4823938221550991   0.9377354660854343   0.7841781755614096   0.9646582786253382   0.29060002806731744   0.3107790311573872   0.7151483918702284   0.5474793189326541   0.7495414433558624   0.711081459141867   0.5262324100657159   0.2743438251430078   0.23349993495091922   0.5984011108937702   0.5431813220599492   0.30366502551638136   0.16228149371853903   0.3459703138347442   0.5581426215688253   0.5986268254939208   0.49529222121125527   0.3194591727307208   0.10592710355255643   0.10480376885873158   0.012898399056156196   0.38172370664528643   0.32174892799114685   0.14014549023339343   0.7222983709888388   0.07094467548789923   0.6066005361209184   0.5926661713007393   0.9727569276329764   0.3598632163460322   0.08036812605520258   0.31832234615773153   0.7392569926820572   0.761462105452262   0.5371868039952534   0.014657320641350158   0.5769754989635182   0.41549179161751776   0.9790441824264281   0.4160304951474294   0.08168327775226286   0.09603261888679697   0.8731170788738717   0.3112267262886978   0.06878487869610667   0.7143089122415105   0.5513681508827248   0.17108123605530437   0.3464865077072679   0.6433642367536113   0.9447676147618065   0.5784150647545651   0.3737295800742915   0.28350102040757913   0.8643994887066039   0.2600927185968336   0.6344725873922343   0.5220389149553172   0.32721268471135045   0.24543539795548341
0.05749708842871614   0.10654712333779937   0.34816850228492235   0.829404902808054   0.9758138106764532   0.010514504451002396   0.4750514234110507   0.5181781765193562   0.9070289319803466   0.29620559220949183   0.9236832725283258   0.3470969404640518   0.5605424242730787   0.6528413554558805   0.9789156577665195   0.7686818757094868   0.1868128441987872   0.36934033504830144   0.11451616905991559   0.5085891571126532   0.5523402568065529   0.8473014200929843   0.7873034843485651   0.2631537591571698   0.4948431683778367   0.7407542967551849   0.43913498206364276   0.4337488563491158   0.5190293577013835   0.7302397923041825   0.9640835586525921   0.9155706798297596   0.6120004257210369   0.4340342000946907   0.04040028612426617   0.5684737393657078   0.05145800144795817   0.7811928446388101   0.061484628357746714   0.799791863656221   0.864645157249171   0.4118525095905087   0.9469684592978311   0.2912027065435678   0.3123049004426181   0.5645510894975244   0.159664974949266   0.028048947386397995   0.8174617320647813   0.8237967927423395   0.7205299928856232   0.5943000910372822   0.2984323743633979   0.093557000438157   0.7564464342330312   0.6787294112075226   0.6864319486423611   0.6595228003434663   0.716046148108765   0.1102556718418149   0.6349739471944029   0.8783299557046562   0.6545615197510183   0.3104638081855939
0.7703287899452319   0.46647744611414754   0.7075930604531872   0.019261101642026112   0.4580238895026138   0.9019263566166231   0.5479280855039211   0.9912121542556281   0.6405621574378324   0.07812956387428363   0.827398092618298   0.39691206321834593   0.3421297830744345   0.9845725634361266   0.07095165838526679   0.7181826520108233   0.6556978344320734   0.32504976309266026   0.3549055102765018   0.6079269801690084   0.02072388723767051   0.44671980738800404   0.7003439905254835   0.2974631719834145   0.2503950972924386   0.9802423612738566   0.9927509300722963   0.2782020703413884   0.7923712077898248   0.07831600465723336   0.4448228445683751   0.28698991608576024   0.15180905035199238   0.00018644078294973408   0.6174247519500772   0.8900778528674144   0.8096792672775579   0.015613877346823103   0.5464730935648103   0.17189520085659107   0.1539814328454845   0.6905641142541629   0.1915675832883086   0.5639682206875827   0.13325754560781397   0.24384430686615877   0.4912235927628251   0.2665050487041682   0.8828624483153754   0.26360194559230227   0.4984726626905288   0.9883029783627798   0.09049124052555056   0.1852859409350689   0.053649818122153685   0.7013130622770196   0.9386821901735581   0.18509950015211918   0.4362250661720765   0.8112352094096053   0.12900292289600027   0.16948562280529605   0.8897519726072661   0.6393400085530142
0.9750214900505157   0.47892150855113325   0.6981843893189575   0.07537178786543147   0.8417639444427019   0.23507720168497448   0.20696079655613242   0.8088667391612633   0.9589014961273264   0.9714752560926723   0.7084881338656036   0.8205637607984835   0.8684102556017759   0.7861893151576033   0.65483831574345   0.11925069852146383   0.9297280654282177   0.6010898150054842   0.2186132495713734   0.3080154891118586   0.8007251425322174   0.4316041922001881   0.3288612769641073   0.6686754805588444   0.8257036524817016   0.9526826836490548   0.6306768876451497   0.593303692693413   0.9839397080389998   0.7176054819640804   0.4237160910890173   0.7844369535321497   0.025038211911673363   0.7461302258714081   0.7152279572234137   0.9638731927336662   0.15662795630989748   0.9599409107138048   0.06038964147996374   0.8446224942122025   0.22689989088167975   0.3588510957083207   0.8417763919085903   0.5366070051003439   0.42617474834946234   0.9272469035081325   0.512915114944483   0.8679315245414995   0.6004710958677607   0.9745642198590777   0.8822382272993333   0.2746278318480865   0.6165313878287608   0.2569587378949974   0.45852213621031607   0.4901908783159368   0.5914931759170875   0.5108285120235893   0.7432941789869024   0.5263176855822705   0.43486521960719005   0.5508876013097844   0.6829045375069387   0.6816951913700681
0.20796532872551027   0.19203650560146374   0.8411281455983484   0.14508818626972425   0.781790580376048   0.26478960209333113   0.32821303065386526   0.27715666172822484   0.18131948450828725   0.2902253822342534   0.4459748033545319   0.0025288298801383765   0.5647880966795265   0.033266644339256024   0.9874526671442158   0.5123379515642016   0.973294920762439   0.5224381323156668   0.2441584881573134   0.986020265981931   0.5384297011552489   0.9715505310058824   0.5612539506503748   0.304325074611863   0.33046437242973864   0.7795140254044186   0.7201258050520264   0.15923688834213873   0.5486737920536907   0.5147244233110875   0.39191277439816113   0.8820802266139139   0.36735430754540344   0.22449904107683405   0.9459379710436292   0.8795513967337755   0.802566210865877   0.19123239673757803   0.9584853038994134   0.36721344516957394   0.8292712901034381   0.6687942644219113   0.7143268157421001   0.38119317918764284   0.29084158894818923   0.6972437334160289   0.15307286509172535   0.07686810457577985   0.9603772165184506   0.9177297080116102   0.43294706003969896   0.9176312162336411   0.41170342446475994   0.4030052847005228   0.04103428564153786   0.035550989619727226   0.04434911691935651   0.17850624362368878   0.09509631459790861   0.15599959288595172   0.2417829060534795   0.9872738468861108   0.13661101069849516   0.7887861477163778
0.4125116159500414   0.31847958246419955   0.4222841949563951   0.40759296852873494   0.12167002700185212   0.6212358490481706   0.2692113298646697   0.3307248639529551   0.1612928104834015   0.7035061410365604   0.8362642698249707   0.413093647719314   0.7495893860186416   0.30050085633603757   0.7952299841834329   0.37754265809958676   0.705240269099285   0.12199461271234881   0.7001336695855243   0.22154306521363504   0.4634573630458056   0.13472076582623804   0.5635226588870291   0.43275691749725725   0.05094574709576421   0.8162411833620385   0.14123846393063402   0.025163948968522296   0.9292757200939121   0.19500533431386785   0.8720271340659643   0.6944390850155672   0.7679829096105106   0.49149919327730746   0.035762864240993536   0.2813454372962532   0.018393523591869028   0.1909983369412699   0.24053288005756066   0.9038027791966665   0.31315325449258397   0.06900372422892109   0.5403992104720363   0.6822597139830314   0.8496958914467784   0.934282958402683   0.9768765515850073   0.24950279648577417   0.7987501443510142   0.11804177504064454   0.8356380876543732   0.2243388475172519   0.8694744242571021   0.9230364407267767   0.963610953588409   0.5298997625016847   0.10149151464659152   0.4315372474494692   0.9278480893474155   0.24855432520543147   0.08309799105472249   0.2405389105081993   0.6873152092898548   0.344751546008765
0.7699447365621385   0.17153518627927822   0.14691599881781842   0.6624918320257336   0.9202488451153601   0.23725222787659517   0.17003944723281114   0.4129890355399594   0.12149870076434591   0.11921045283595064   0.3344013595784379   0.1886501880227075   0.2520242765072438   0.19617401210917396   0.37079040599002894   0.6587504255210228   0.1505327618606523   0.7646367646597048   0.4429423166426135   0.41019610031559134   0.06743477080592979   0.5240978541515054   0.7556271073527587   0.06544455430682636   0.2974900342437913   0.3525626678722272   0.6087111085349404   0.4029527222810928   0.3772411891284312   0.11531043999563202   0.4386716613021292   0.9899636867411334   0.25574248836408525   0.9960999871596814   0.1042703017236913   0.8013134987184258   0.0037182118568414753   0.7999259750505074   0.7334798957336623   0.14256307319740305   0.8531854499961892   0.0352892103908027   0.2905375790910488   0.7323669728818117   0.7857506791902594   0.5111913562392972   0.5349104717382901   0.6669224185749854   0.48826064494646815   0.1586286883670701   0.9261993632033497   0.26396969629389255   0.11101945581803696   0.04331824837143805   0.4875277019012205   0.27400600955275917   0.8552769674539517   0.047218261211756665   0.38325740017752924   0.4726925108343333   0.8515587555971103   0.24729228616124924   0.6497775044438668   0.33012943763693026
0.998373305600921   0.21200307577044653   0.35923992535281807   0.5977624647551185   0.2126226264106616   0.7008117195311493   0.8243294536145279   0.9308400461801332   0.7243619814641935   0.5421830311640792   0.8981300904111782   0.6668703498862406   0.6133425256461565   0.4988647827926411   0.4106023885099577   0.39286434033348144   0.7580655581922048   0.4516465215808845   0.02734498833242849   0.9201718294991481   0.9065068025950946   0.20435423541963524   0.3775674838885616   0.590042391862218   0.9081334969941736   0.9923511596491887   0.018327558535743575   0.9922799271070993   0.695510870583512   0.29153944011803945   0.1939981049212156   0.061439880926966194   0.9711488891193185   0.7493564089539603   0.29586801451003736   0.39456953104072556   0.357806363473162   0.25049162616131915   0.8852656260000796   0.001705190707244134   0.5997408052809572   0.7988451045804347   0.8579206376676511   0.08153336120809598   0.6932340026858625   0.5944908691607994   0.48035315377908955   0.4914909693458781   0.785100505691689   0.6021397095116108   0.46202559524334597   0.4992110422387787   0.08958963510817698   0.3106002693935713   0.26802749032213036   0.43777116131181254   0.11844074598885847   0.561243860439611   0.9721594758120929   0.04320163027108694   0.7606343825156965   0.3107522342782919   0.08689384981201334   0.04149643956384281
0.1608935772347393   0.5119071296978572   0.22897321214436217   0.9599630783557468   0.46765957454887674   0.9174162605370577   0.7486200583652727   0.46847210900986874   0.6825590688571878   0.315276551025447   0.28659446312192666   0.96926106677109   0.5929694337490108   0.004676281631875707   0.018566972799796317   0.5314899054592775   0.4745286877601523   0.44343242119226467   0.04640749698770332   0.48828827518819057   0.7138943052444559   0.1326801869139728   0.95951364717569   0.44679183562434777   0.5530007280097166   0.6207730572161155   0.7305404350313278   0.4868287572686009   0.08534115346083981   0.7033567966790578   0.9819203766660551   0.01835664825873221   0.40278208460365206   0.3880802456536108   0.6953259135441284   0.04909558148764218   0.8098126508546413   0.3834039640217351   0.6767589407443322   0.5176056760283647   0.335283963094489   0.9399715428294705   0.6303514437566289   0.029317400840174097   0.6213896578500332   0.8072913559154976   0.6708377965809389   0.5825255652158263   0.06838892984031661   0.18651829869938208   0.9402973615496111   0.09569680794722539   0.9830477763794768   0.48316150202032426   0.9583769848835559   0.07734015968849318   0.5802656917758248   0.09508125636671343   0.26305107133942746   0.028244578200851   0.7704530409211835   0.7116772923449783   0.5862921305950952   0.5106389021724863
0.4351690778266945   0.7717057495155079   0.9559406868384664   0.4813215013323122   0.8137794199766614   0.9644143936000102   0.28510289025752755   0.8987959361164859   0.7453904901363447   0.7778960949006282   0.3448055287079165   0.8030991281692605   0.7623427137568679   0.2947345928803039   0.3864285438243606   0.7257589684807674   0.1820770219810432   0.1996533365135905   0.12337747248493316   0.6975143902799164   0.4116239810598597   0.4879760441686122   0.5370853418898379   0.18687548810743   0.9764549032331652   0.7162702946531043   0.5811446550513715   0.7055539867751177   0.1626754832565039   0.7518559010530941   0.2960417647938439   0.8067580506586318   0.4172849931201592   0.9739598061524659   0.9512362360859274   0.0036589224893713653   0.6549422793632913   0.6792252132721619   0.5648076922615668   0.27789995400860407   0.47286525738224805   0.47957187675857144   0.44143021977663366   0.5803855637286877   0.06124127632238835   0.9915958325899593   0.9043448778867957   0.3935100756212577   0.0847863730892231   0.275325537936855   0.32320022283542427   0.6879560888461399   0.9221108898327192   0.523469636883761   0.027158458041580392   0.8811980381875081   0.5048258967125601   0.5495098307312951   0.075922221955653   0.8775391156981367   0.8498836173492688   0.8702846174591331   0.5111145296940862   0.5996391616895327
0.3770183599670207   0.39071274070056167   0.06968430991745254   0.019253597960844956   0.31577708364463236   0.3991169081106024   0.1653394320306568   0.6257435223395873   0.23099071055540923   0.12379137017374738   0.8421392091952324   0.9377874334934473   0.30887982072269005   0.6003217332899864   0.8149807511536521   0.056589395305939226   0.80405392401013   0.05081190255869131   0.7390585291979991   0.1790502796078025   0.9541703066608612   0.18052728509955818   0.22794399950391292   0.5794111179182698   0.5771519466938406   0.7898145443989965   0.1582596895864604   0.5601575199574249   0.26137486304920826   0.3906976362883941   0.9929202575558036   0.9344139976178376   0.030384152493799013   0.26690626611464674   0.1507810483605711   0.9966265641243903   0.721504331771109   0.6665845328246603   0.335800297206919   0.9400371688184511   0.917450407760979   0.6157726302659691   0.5967417680089199   0.7609868892106486   0.9632801011001176   0.4352453451664109   0.36879776850500695   0.18157577129237876   0.38612815440627707   0.6454308007674143   0.21053807891854656   0.6214182513349539   0.12475329135706884   0.2547331644790203   0.21761782136274296   0.6870042537171163   0.09436913886326982   0.9878268983643735   0.06683677300217188   0.6903776895927258   0.37286480709216085   0.3212423655397132   0.7310364757952529   0.7503405207742747
0.4554143993311819   0.7054697352737441   0.13429470778633298   0.9893536315636262   0.49213429823106425   0.2702243901073333   0.765496939281326   0.8077778602712474   0.10600614382478714   0.6247935893399189   0.5549588603627794   0.18635960893629352   0.9812528524677183   0.37006042486089863   0.3373410390000365   0.4993553552191773   0.8868837136044485   0.3822335264965251   0.2705042659978646   0.8089776656264515   0.5140189065122877   0.06099116095681192   0.5394677902026117   0.058637144852176665   0.058604507181105756   0.35552142568306777   0.40517308241627875   0.06928351328855051   0.5664702089500415   0.08529703557573445   0.6396761431349527   0.2615056530173031   0.4604640651252544   0.4605034462358155   0.08471728277217325   0.07514604408100957   0.4792112126575361   0.09044302137491689   0.7473762437721367   0.5757906888618323   0.5923274990530876   0.7082094948783918   0.47687197777427215   0.7668130232353808   0.07830859254079992   0.6472183339215799   0.9374041875716604   0.7081758783832042   0.019704085359694163   0.29169690823851213   0.5322311051553816   0.6388923650946536   0.4532338764096526   0.20639987266277765   0.8925549620204289   0.3773867120773506   0.9927698112843982   0.7458964264269621   0.8078376792482557   0.30224066799634103   0.5135585986268622   0.6554534050520452   0.060461435476118944   0.7264499791345087
0.9212310995737746   0.9472439101736535   0.5835894577018468   0.9596369558991279   0.8429225070329747   0.3000255762520736   0.6461852701301863   0.2514610775159237   0.8232184216732805   0.00832866801356149   0.11395416497480469   0.61256871242127   0.3699845452636279   0.8019287953507839   0.22139920295437573   0.23518200034391945   0.37721473397922967   0.05603236892382171   0.41356152370612004   0.9329413323475785   0.8636561353523674   0.4005789638717765   0.35310008823000105   0.20649135321306972   0.9424250357785928   0.453335053698123   0.7695106305281543   0.24685439731394182   0.09950252874561814   0.15330947744604942   0.12332536039796792   0.9953933197980182   0.27628410707233764   0.14498080943248792   0.00937119542316323   0.3828246073767481   0.9062995618087097   0.3430520140817041   0.7879719924687875   0.14764260703282867   0.5290848278294801   0.28701964515788236   0.3744104687626675   0.21470127468525022   0.6654286924771127   0.8864406812861059   0.0213103805326664   0.008209921472180517   0.7230036566985198   0.4331056275879829   0.2517997500045121   0.7613555241582387   0.6235011279529017   0.2797961501419335   0.1284743896065442   0.7659622043602206   0.347217020880564   0.13481534070944554   0.11910319418338096   0.3831375969834725   0.4409174590718543   0.7917633266277414   0.3311312017145935   0.2354949899506438
0.9118326312423742   0.504743681469859   0.956720732951926   0.02079371526539358   0.24640393876526157   0.6183030001837532   0.9354103524192596   0.012583793793213062   0.5234002820667417   0.18519737259577027   0.6836106024147475   0.25122826963497435   0.8998991541138401   0.9054012224538368   0.5551362128082032   0.4852660652747538   0.5526821332332761   0.7705858817443912   0.43603301862482235   0.10212846829128133   0.11176467416142181   0.9788225551166498   0.10490181691022887   0.8666334783406375   0.19993204291904762   0.47407887364679074   0.1481810839583029   0.8458397630752439   0.9535281041537861   0.8557758734630376   0.21277073153904333   0.8332559692820308   0.43012782208704425   0.6705785008672673   0.5291601291242959   0.5820276996470565   0.5302286679732041   0.7651772784134305   0.9740239163160925   0.09676163437230272   0.977546534739928   0.9945913966690393   0.5379908976912703   0.9946331660810214   0.8657818605785063   0.0157688415523895   0.43308908078104136   0.12799968774038387   0.6658498176594586   0.5416899679055988   0.2849079968227385   0.2821599246651399   0.7123217135056725   0.6859140944425611   0.07213726528369514   0.44890395538310907   0.28219389141862833   0.015335593575293849   0.5429771361593992   0.8668762557360525   0.7519652234454242   0.2501583151618633   0.5689532198433067   0.7701146213637499
0.7744186887054961   0.255566918492824   0.03096232215203648   0.7754814552827284   0.9086368281269899   0.2397980769404345   0.5978732413709951   0.6474817675423445   0.24278701046753126   0.6981081090348358   0.31296524454825664   0.36532184287720465   0.5304652969618586   0.012194014592274566   0.2408279792645615   0.9164178874940956   0.24827140554323035   0.9968584210169807   0.6978508431051622   0.04954163175804307   0.4963061820978062   0.7467001058551174   0.1288976232618555   0.27942701039429324   0.7218874933923101   0.4911331873622934   0.097935301109819   0.5039455551115648   0.8132506652653202   0.2513351104218589   0.5000620597388239   0.8564637875692203   0.5704636547977889   0.5532270013870232   0.18709681519056723   0.4911419446920156   0.039998357835930295   0.5410329867947485   0.9462688359260057   0.5747240571979201   0.7917269522927   0.5441745657777679   0.24841799282084354   0.5251824254398769   0.2954207701948937   0.7974744599226504   0.11952036955898804   0.2457554150455837   0.5735332768025836   0.30634127256035704   0.021585068449169038   0.7418098599340189   0.7602826115372634   0.05500616213849816   0.5215230087103452   0.8853460723647986   0.18981895673947444   0.501779160751475   0.3344261935197779   0.394204127672783   0.14982059890354416   0.9607461739567265   0.3881573575937722   0.8194800704748629
0.3580936466108442   0.41657160817895855   0.13973936477292864   0.294297645034986   0.0626728764159505   0.6190971482563081   0.020218995213940612   0.048542229989402275   0.48913959961336684   0.31275587569595104   0.9986339267647716   0.3067323700553834   0.7288569880761034   0.25774971355745285   0.4771109180544264   0.4213862976905848   0.539038031336629   0.7559705528059779   0.1426847245346485   0.027182170017801797   0.3892174324330848   0.7952243788492515   0.7545273669408763   0.20770209954293883   0.03112378582224062   0.3786527706702929   0.6147880021679477   0.9134044545079528   0.9684509094062901   0.7595556224139848   0.594569006954007   0.8648622245185505   0.47931130979292325   0.4467997467180338   0.5959350801892355   0.5581298544631672   0.7504543217168198   0.18905003316058092   0.11882416213480906   0.1367435567725824   0.21141629038019083   0.4330794803546031   0.9761394376001605   0.10956138675478061   0.822198857947106   0.6378551015053516   0.22161207065928423   0.9018592872118417   0.7910750721248654   0.2592023308350587   0.6068240684913365   0.9884548327038889   0.8226241627185752   0.4996467084210739   0.012255061537329498   0.12359260818533833   0.34331285292565195   0.0528469617030401   0.416319981348094   0.5654627537221711   0.5928585312088321   0.8637969285424592   0.29749581921328494   0.4287191969495887
0.3814422408286413   0.4307174481878561   0.3213563816131244   0.3191578101948081   0.5592433828815353   0.7928623466825045   0.09974431095384016   0.4172985229829663   0.7681683107566699   0.5336600158474458   0.4929202424625036   0.4288436902790774   0.9455441480380947   0.03401330742637191   0.48066518092517413   0.3052510820937391   0.6022312951124428   0.9811663457233318   0.0643451995770801   0.7397883283715679   0.0093727639036106   0.11736941718087263   0.7668493803637951   0.31106913142197923   0.6279305230749693   0.6866519689930165   0.4454929987506707   0.9919113212271711   0.06868714019343396   0.893789622310512   0.3457486877968306   0.5746127982442047   0.300518829436764   0.3601296064630662   0.852828445334327   0.14576910796512735   0.3549746813986693   0.32611629903669426   0.37216326440915287   0.8405180258713882   0.7527433862862265   0.3449499533133625   0.30781806483207275   0.10072969749982028   0.743370622382616   0.22758053613248985   0.5409686844682776   0.7896605660778411   0.11544009930764665   0.5409285671394733   0.09547568571760687   0.7977492448506699   0.04675295911421269   0.6471389448289614   0.7497269979207762   0.22313644660646512   0.7462341296774487   0.28700933836589515   0.8968985525864493   0.07736733864133778   0.3912594482787794   0.9608930393292009   0.5247352881772964   0.23684931276994953
0.6385160619925528   0.6159430860158384   0.2169172233452237   0.13611961527012925   0.895145439609937   0.38836254988334856   0.6759485388769461   0.3464590491922882   0.7797053403022903   0.8474339827438752   0.5804728531593393   0.5487098043416183   0.7329523811880776   0.20029503791491382   0.8307458552385629   0.32557335773515317   0.9867182515106289   0.9132856995490186   0.9338473026521136   0.2482060190938154   0.5954588032318495   0.9523926602198177   0.40911201447481715   0.01135670632386586   0.9569427412392967   0.33644957420397936   0.19219479112959348   0.8752370910537366   0.061797301629359674   0.9480870243206309   0.5162462522526474   0.5287780418614484   0.2820919613270694   0.10065304157675561   0.9357733990933081   0.9800682375198301   0.5491395801389918   0.9003580036618418   0.10502754385474522   0.6544948797846769   0.5624213286283628   0.9870723041128231   0.1711802412026316   0.4062888606908615   0.9669625253965134   0.03467964389300537   0.7620682267278144   0.39493215436699564   0.010019784157216716   0.698230069689026   0.569873435598221   0.519695063313259   0.948222482527857   0.7501430453683952   0.05362718334557358   0.9909170214518106   0.6661305212007876   0.6494900037916396   0.11785378425226542   0.01084878393198058   0.1169909410617959   0.7491320001297977   0.012826240397520193   0.35635390414730367
0.5545696124334331   0.7620596960169747   0.8416459991948886   0.9500650434564422   0.5876070870369197   0.7273800521239693   0.07957777246707416   0.5551328890894466   0.577587302879703   0.02914998243494328   0.5097043368688532   0.03543782577618752   0.6293648203518459   0.2790069370665481   0.45607715352327965   0.04452080432437687   0.9632342991510583   0.6295169332749085   0.3382233692710142   0.033672020392396286   0.8462433580892624   0.8803849331451107   0.32539712887349403   0.6773181162450926   0.2916737456558293   0.11832523712813607   0.48375112967860545   0.7272530727886504   0.7040666586189096   0.3909451850041668   0.40417335721153125   0.17212018369920384   0.12647935573920663   0.3617952025692235   0.8944690203426781   0.13668235792301633   0.49711453538736067   0.08278826550267543   0.4383918668193984   0.09216155359863946   0.5338802362363023   0.4532713322277669   0.10016849754838421   0.05848953320624318   0.68763687814704   0.5728863990826562   0.7747713686748902   0.3811714169611506   0.3959631324912106   0.4545611619545201   0.29102023899628476   0.6539183441725002   0.691896473872301   0.06361597695035331   0.8868468817847535   0.4817981604732963   0.5654171181330944   0.7018207743811298   0.9923778614420754   0.34511580255027996   0.06830258274573374   0.6190325088784544   0.5539859946226771   0.2529542489516405
0.5344223465094313   0.16576117665068746   0.4538174970742928   0.19446471574539734   0.8467854683623914   0.5928747775680313   0.6790461283994026   0.8132932987842467   0.45082233587118076   0.1383136156135112   0.3880258894031179   0.15937495461174658   0.7589258619988797   0.07469763866315787   0.5011790076183644   0.6775767941384503   0.19350874386578532   0.3728768642820281   0.5088011461762889   0.3324609915881703   0.1252061611200516   0.7538443554035736   0.954815151553612   0.07950674263652979   0.5907838146106202   0.5880831787528862   0.5009976544793191   0.8850420268911324   0.7439983462482288   0.995208401184855   0.8219515260799165   0.0717487281068857   0.29317601037704805   0.8568947855713438   0.4339256366767986   0.9123737734951392   0.5342501483781683   0.7821971469081859   0.9327466290584342   0.23479697935668886   0.340741404512383   0.4093202826261578   0.4239454828821453   0.9023359877685185   0.21553524339233143   0.6554759272225841   0.4691303313285333   0.8228292451319887   0.6247514287817112   0.06739274846969788   0.9681326768492142   0.9377872182408563   0.8807530825334824   0.07218434728484295   0.14618115076929766   0.8660384901339706   0.5875770721564344   0.2152895617134992   0.712255514092499   0.9536647166388315   0.05332692377826602   0.4330924148053133   0.7795088850340648   0.7188677372821426
0.712585519265883   0.023772132179155494   0.35556340215191956   0.8165317495136241   0.49705027587355155   0.3682962049565714   0.8864330708233862   0.9937025043816353   0.8722988470918404   0.3009034564868735   0.9183003939741721   0.05591528614077899   0.991545764558358   0.22871910920203056   0.7721192432048744   0.18987679600680837   0.40396869240192357   0.013429547488531361   0.05986372911237536   0.2362120793679769   0.35064176862365753   0.5803371326832181   0.28035484407831057   0.5173443420858342   0.6380562493577746   0.5565650005040625   0.9247914419263911   0.7008125925722102   0.14100597348422297   0.18826879554749118   0.038358371103004794   0.7071100881905749   0.26870712639238264   0.8873653390606177   0.12005797712883273   0.651194802049796   0.27716136183402473   0.6586462298585871   0.34793873392395835   0.4613180060429875   0.8731926694321012   0.6452166823700558   0.288075004811583   0.22510592667501064   0.5225509008084436   0.06487954968683772   0.007720160733272416   0.7077615845891764   0.884494651450669   0.5083145491827752   0.0829287188068814   0.006948992016966175   0.743488677966446   0.320045753635284   0.044570347703876606   0.2998389038263913   0.4747815515740634   0.43268041457466627   0.9245123705750439   0.6486441017765954   0.19762018974003867   0.7740341847160792   0.5765736366510855   0.18732609573360784
0.32442752030793753   0.12881750234602338   0.2884986318395026   0.9622201690585972   0.801876619499494   0.06393795265918566   0.28077847110623017   0.2544585844694208   0.917381968048825   0.5556234034764105   0.19784975229934876   0.24750959245245466   0.17389329008237894   0.23557764984112653   0.15327940459547215   0.9476706886260634   0.6991117385083155   0.8028972352664602   0.22876703402042828   0.29902658684946803   0.5014915487682768   0.028863050550381072   0.6521933973693428   0.11170049111586017   0.17706402846033933   0.9000455482043577   0.3636947655298402   0.14948032205726294   0.37518740896084535   0.836107595545172   0.08291629442361004   0.8950217375878421   0.45780544091202036   0.2804841920687615   0.8850665421242613   0.6475121451353875   0.28391215082964144   0.044906542227635   0.7317871375287891   0.6998414565093241   0.5848004123213258   0.24200930696117476   0.5030201035083609   0.4008148696598561   0.08330886355304896   0.2131462564107937   0.8508267061390181   0.2891143785439959   0.9062448350927096   0.313100708206436   0.48713194060917797   0.13963405648673294   0.5310574261318642   0.476993112661264   0.40421564618556793   0.24461231889889082   0.07325198521984388   0.19650892059250247   0.5191491040613067   0.5971001737635033   0.7893398343902025   0.15160237836486745   0.7873619665325174   0.8972587172541793
0.2045394220688766   0.9095930714036927   0.2843418630241566   0.49644384759432325   0.12123055851582765   0.696446814992899   0.4335151568851385   0.20732946905032737   0.21498572342311803   0.38334610678646297   0.9463832162759604   0.06769541256359443   0.6839282972912538   0.906352994125199   0.5421675700903925   0.8230830936647037   0.6106763120714099   0.7098440735326965   0.023018466029085912   0.22598291990120023   0.8213364776812074   0.5582416951678291   0.23565649949656842   0.32872420264702096   0.6167970556123308   0.6486486237641363   0.9513146364724118   0.8322803550526977   0.4955664970965032   0.9522018087712374   0.5177994795872733   0.6249508860023703   0.28058077367338513   0.5688557019847744   0.5714162633113129   0.5572554734387759   0.5966524763821314   0.6625027078595754   0.02924869322092029   0.7341723797740722   0.9859761643107215   0.9526586343268789   0.006230227191834381   0.508189459872872   0.1646396866295141   0.3944169391590498   0.770573727695266   0.17946525722585108   0.5478426310171832   0.7457683153949134   0.8192590912228541   0.3471849021731534   0.05227613392068009   0.793566506623676   0.3014596116355808   0.7222340161707831   0.7716953602472949   0.22471080463890158   0.730043348324268   0.16497854273200724   0.17504288386516356   0.5622080967793261   0.7007946551033477   0.43080616295793495
0.18906671955444204   0.6095494624524473   0.6945644279115133   0.9226167030850629   0.02442703292492796   0.21513252329339755   0.9239907002162473   0.7431514458592119   0.4765844019077447   0.46936420789848415   0.10473160899339316   0.39596654368605844   0.4243082679870646   0.6757977012748081   0.8032719973578124   0.6737325275152753   0.6526129077397697   0.45108689663590656   0.07322864903354438   0.5087539847832682   0.4775700238746061   0.8888787998565804   0.3724339939301967   0.07794782182533318   0.2885033043201641   0.279329337404133   0.6778695660186834   0.15533111874027022   0.2640762713952361   0.0641968141107355   0.7538788658024361   0.41217967288105833   0.7874918694874914   0.5948326062122513   0.649147256809043   0.016213129194999888   0.36318360150042683   0.9190349049374432   0.8458752594512305   0.3424806016797245   0.7105706937606572   0.46794800830153666   0.7726466104176862   0.8337266168964563   0.23300066988605106   0.5790692084449562   0.40021261648748946   0.7557787950711232   0.944497365565887   0.2997398710408232   0.7223430504688061   0.6004476763308529   0.6804210941706509   0.23554305693008776   0.96846418466637   0.18826800344979464   0.8929292246831595   0.6407104507178364   0.319316927857327   0.17205487425479474   0.5297456231827327   0.7216755457803932   0.47344166840609647   0.8295742725750702
0.8191749294220755   0.2537275374788565   0.7007950579884102   0.9958476556786139   0.5861742595360244   0.6746583290339002   0.3005824415009208   0.24006886060749064   0.6416768939701375   0.374918457993077   0.5782393910321147   0.6396211842766376   0.9612557997994866   0.13937540106298923   0.6097752063657448   0.451353180826843   0.06832657511632709   0.49866495034515285   0.29045827850841777   0.2792983065720483   0.5385809519335945   0.7769894045647596   0.8170166101023213   0.449724033996978   0.7194060225115189   0.5232618670859032   0.11622155211391101   0.4538763783183642   0.13323176297549447   0.8486035380520028   0.8156391106129902   0.21380751771087356   0.491554869005357   0.47368508005892584   0.23739971958087547   0.5741863334342359   0.5302990692058704   0.3343096789959366   0.6276245132151307   0.12283315260739289   0.4619724940895434   0.8356447286507838   0.337166234706713   0.8435348460353446   0.923391542155949   0.05865532408602411   0.5201496246043917   0.3938108120383666   0.20398551964443004   0.535393457000121   0.4039280724904807   0.9399344337200024   0.07075375666893557   0.6867899189481181   0.5882889618774905   0.7261269160091288   0.5791988876635785   0.2131048388891923   0.35088924229661494   0.1519405825748929   0.048899818457708126   0.8787951598932556   0.7232647290814843   0.029107429967500015
0.5869273243681647   0.0431504312424719   0.3860984943747713   0.1855725839321554   0.6635357822122159   0.9844951071564478   0.8659488697703797   0.7917617718937888   0.4595502625677858   0.4491016501563268   0.4620207972798989   0.8518273381737864   0.38879650589885023   0.7623117312082086   0.8737318354024085   0.12570042216465765   0.8095976182352717   0.5492068923190163   0.5228425931057935   0.9737598395897648   0.7606977997775635   0.6704117324257607   0.7995778640243093   0.9446524096222647   0.17377047540939874   0.6272613011832888   0.41347936964953796   0.7590798256901093   0.510234693197183   0.642766194026841   0.5475304998791584   0.9673180537963205   0.050684430629397134   0.1936645438705142   0.0855097025992594   0.11549071562253405   0.6618879247305469   0.4313528126623056   0.2117778671968509   0.9897902934578764   0.8522903064952753   0.8821459203432892   0.6889352740910574   0.01603045386811166   0.0915925067177118   0.21173418791752854   0.8893574100667481   0.07137804424584693   0.9178220313083131   0.5844728867342398   0.47587804041721016   0.3122982185557376   0.4075873381111301   0.9417066927073987   0.9283475405380518   0.3449801647594171   0.356902907481733   0.7480421488368846   0.8428378379387924   0.22948944913688304   0.6950149827511861   0.31668933617457895   0.6310599707419415   0.23969915567900665
0.8427246762559107   0.43454341583128975   0.9421246966508842   0.223668701810895   0.751132169538199   0.22280922791376118   0.05276728658413603   0.15229065756504806   0.8333101382298859   0.6383363411795214   0.5768892461669258   0.8399924390093104   0.4257228001187558   0.6966296484721227   0.648541705628874   0.49501227424989336   0.06881989263702279   0.9485874996352381   0.8057038676900816   0.2655228251130103   0.3738049098858367   0.6318981634606592   0.1746438969481401   0.025823669434003656   0.531080233629926   0.19735474762936947   0.23251920029725595   0.8021549676231087   0.779948064091727   0.9745455197156083   0.1797519137131199   0.6498643100580606   0.946637925861841   0.33620917853608684   0.602862667546194   0.8098718710487501   0.5209151257430853   0.6395795300639642   0.95432096191732   0.3148595967988568   0.4520952331060625   0.690992030428726   0.14861709422723837   0.04933677168584649   0.07829032322022578   0.059093866968066816   0.9739731972790983   0.023513102251842836   0.5472100895902998   0.8617391193386973   0.7414539969818423   0.22135813462873416   0.7672620254985728   0.8871935996230891   0.5617020832687224   0.5714938245706735   0.8206240996367318   0.5509844210870022   0.9588394157225284   0.7616219535219234   0.2997089738936465   0.911404891023038   0.00451845380520837   0.4467623567230666
0.847613740787584   0.220412860594312   0.85590135957797   0.3974255850372201   0.7693234175673582   0.1613189936262452   0.8819281622988717   0.37391248278537725   0.2221133279770584   0.29957987428754784   0.1404741653170294   0.1525543481566431   0.45485130247848554   0.4123862746644588   0.578772082048307   0.5810605235859695   0.6342272028417538   0.8614018535774566   0.6199326663257786   0.8194385700640462   0.33451822894810734   0.9499969625544186   0.6154142125205703   0.37267621334097956   0.48690448816052334   0.7295841019601066   0.7595128529426003   0.9752506283037594   0.7175810705931651   0.5682651083338613   0.8775846906437286   0.6013381455183822   0.49546774261610677   0.2686852340463135   0.7371105253266992   0.44878379736173907   0.04061644013762117   0.8562989593818547   0.15833844327839217   0.8677232737757695   0.40638923729586734   0.994897105804398   0.5384057769526136   0.04828470371172339   0.07187100834776003   0.04490014324997955   0.9229915644320433   0.6756084903707439   0.5849665201872367   0.315316041289873   0.16347871148944307   0.7003578620669844   0.8673854495940716   0.7470509329560117   0.2858940208457146   0.09901971654860223   0.37191770697796483   0.47836569890969816   0.5487834955190154   0.6502359191868632   0.33130126684034367   0.6220667395278434   0.39044505224062326   0.7825126454110937
0.9249120295444763   0.6271696337234454   0.8520392752880097   0.7342279416993702   0.8530410211967162   0.5822694904734658   0.9290477108559664   0.05861945132862639   0.26807450100947955   0.2669534491835928   0.7655689993665233   0.358261589261642   0.400689051415408   0.5199025162275811   0.47967497852080876   0.2592418727130398   0.028771344437443204   0.04153681731788299   0.9308914830017934   0.6090059535261766   0.6974700775970996   0.41947007779003953   0.54044643076117   0.826493308115083   0.7725580480526233   0.7923004440665942   0.6884071554731603   0.09226536641571279   0.9195170268559071   0.21003095359312837   0.759359444617194   0.03364591508708639   0.6514425258464275   0.9430775044095355   0.9937904452506706   0.6753843258254444   0.2507534744310195   0.4231749881819544   0.514115466729862   0.4161424531124046   0.22198212999357625   0.3816381708640714   0.5832239837280686   0.807136499586228   0.5245120523964767   0.9621680930740318   0.04277755296689855   0.980643191471145   0.7519540043438534   0.16986764900743773   0.3543703974937382   0.8883778250554322   0.8324369774879464   0.9598366954143094   0.5950109528765443   0.8547319099683458   0.1809944516415189   0.0167591910047738   0.6012205076258735   0.17934758414290142   0.9302409772104995   0.5935842028228194   0.08710504089601163   0.7632051310304968
0.7082588472169232   0.21194603195874798   0.5038810571679431   0.9560686314442688   0.18374679482044648   0.24977793888471608   0.46110350420104446   0.9754254399731238   0.4317927904765931   0.07991028987727836   0.10673310670730628   0.08704761491769164   0.5993558129886467   0.120073594462969   0.511722153830762   0.23231570494934584   0.4183613613471278   0.1033144034581952   0.9105016462048885   0.05296812080644443   0.48812038413662834   0.5097302006353758   0.8233966053088768   0.28976298977594767   0.7798615369197052   0.2977841686766278   0.31951554814093386   0.3336943583316789   0.5961147420992587   0.04800622979191176   0.8584120439398893   0.358268918358555   0.16432195162266564   0.9680959399146334   0.751678937232583   0.27122130344086337   0.5649661386340189   0.8480223454516644   0.23995678340182106   0.038905598491517555   0.14660477728689117   0.7447079419934692   0.32945513719693253   0.9859374776850731   0.6584843931502627   0.23497774135809338   0.5060585318880557   0.6961744879091255   0.8786228562305576   0.9371935726814655   0.18654298374712186   0.36248012957744663   0.2825081141312989   0.8891873428895538   0.3281309398072325   0.004211211218891605   0.11818616250863326   0.9210914029749203   0.5764520025746495   0.7329899077780282   0.5532200238746143   0.07306905752325597   0.3364952191728284   0.6940843092865107
0.40661524658772313   0.3283611155297868   0.007040081975895824   0.7081468316014375   0.7481308534374603   0.09338337417169341   0.5009815500878402   0.011972343692312055   0.8695079972069027   0.15618980149022788   0.31443856634071826   0.6494922141148655   0.5869998830756038   0.2670024586006741   0.9863076265334857   0.6452810028959738   0.46881372056697057   0.34591105562575375   0.4098556239588363   0.9122910951179456   0.9155936966923562   0.27284199810249776   0.07336040478600793   0.21820678583143494   0.5089784501046332   0.944480882572711   0.0663203228101121   0.5100599542299974   0.7608475966671728   0.8510975084010176   0.565338772722272   0.49808761053768535   0.8913395994602701   0.6949077069107897   0.25090020638155375   0.8485953964228199   0.3043397163846662   0.42790524831011556   0.264592579848068   0.2033143935268461   0.8355259958176956   0.08199419268436182   0.8547369558892317   0.2910232984089005   0.9199322991253394   0.809152194581864   0.7813765511032238   0.07281651257746556   0.4109538490207062   0.864671312009153   0.7150562282931117   0.5627565583474682   0.6501062523535334   0.013573803608135458   0.14971745557083965   0.06466894780978279   0.7587666528932634   0.31866609669734575   0.898817249189286   0.21607355138696285   0.4544269365085971   0.8907608483872301   0.6342246693412179   0.01275915786011674
0.6189009406909015   0.8087666557028683   0.7794877134519862   0.7217358594512162   0.6989686415655622   0.9996144611210043   0.9981111623487625   0.6489193468737506   0.288014792544856   0.13494314911185123   0.28305493405565085   0.08616278852628254   0.6379085401913226   0.12136934550371578   0.1333374784848112   0.021493840716499752   0.8791418872980593   0.80270324880637   0.23452022929552527   0.8054202893295369   0.42471495078946214   0.9119424004191399   0.6002955599543074   0.7926611314694202   0.8058140100985606   0.10317574471627153   0.8208078465023211   0.07092527201820392   0.10684536853299843   0.10356128359526723   0.8226966841535586   0.42200592514445323   0.8188305759881425   0.9686181344834159   0.5396417500979077   0.3358431366181707   0.18092203579681984   0.8472487889797002   0.40630427161309657   0.314349295901671   0.3017801484987606   0.04454554017333017   0.1717840423175713   0.508929006572134   0.8770651977092985   0.1326031397541903   0.571488482363264   0.716267875102714   0.07125118761073784   0.029427395037918785   0.7506806358609428   0.64534260308451   0.9644058190777394   0.9258661114426515   0.9279839517073842   0.22333667794005674   0.14557524308959696   0.9572479769592356   0.38834220160947647   0.8874935413218861   0.9646532072927771   0.10999918797953537   0.9820379299963798   0.573144245420215
0.6628730587940165   0.06545364780620519   0.8102538876788086   0.06421523884808099   0.785807861084718   0.9328505080520149   0.23876540531554466   0.3479473637453671   0.7145566734739802   0.9034231130140961   0.48808476945460183   0.7026047606608571   0.7501508543962409   0.9775570015714445   0.5601008177472175   0.4792680827208004   0.6045756113066438   0.02030902461220898   0.17175861613774113   0.5917745413989144   0.6399224040138668   0.9103098366326736   0.18972068614136123   0.018630295978699314   0.9770493452198502   0.8448561888264684   0.3794667984625526   0.9544150571306184   0.19124148413513217   0.9120056807744535   0.14070139314700797   0.6064676933852512   0.476684810661152   0.008582567760357436   0.6526166236924061   0.9038629327243941   0.7265339562649111   0.03102556618891289   0.09251580594518859   0.42459485000359376   0.12195834495826728   0.01071654157670391   0.9207571898074475   0.8328203086046794   0.48203594094440055   0.1004067049440303   0.7310365036660863   0.81419001262598   0.5049865957245503   0.25555051611756185   0.35156970520353364   0.8597749554953618   0.3137451115894181   0.3435448353431083   0.21086831205652565   0.2533072621101105   0.8370603009282661   0.3349622675827509   0.5582516883641194   0.3494443293857164   0.11052634466335502   0.303936701393838   0.4657358824189309   0.9248494793821227
0.9885679997050877   0.2932201598171341   0.5449786926114835   0.09202917077744328   0.5065320587606872   0.1928134548731038   0.8139421889453972   0.27783915815146326   0.0015454630361369113   0.9372629387555419   0.4623724837418635   0.4180642026561015   0.6878003514467188   0.5937181034124336   0.2515041716853379   0.164756940545991   0.8507400505184526   0.2587558358296827   0.6932524833212184   0.8153126111602746   0.7402137058550976   0.9548191344358447   0.2275166009022875   0.890463131778152   0.7516457061500099   0.6615989746187106   0.6825379082908041   0.7984339610007087   0.24511364738932268   0.4687855197456068   0.8685957193454069   0.5205948028492454   0.24356818435318575   0.5315225809900649   0.4062232356035434   0.10253060019314394   0.5557678329064669   0.9378044775776313   0.15471906391820556   0.937773659647153   0.7050277823880143   0.6790486417479485   0.46146658059698714   0.12246104848687832   0.9648140765329167   0.7242295073121039   0.23394997969469963   0.23199791670872635   0.21316837038290684   0.06263053269339328   0.5514120714038956   0.43356395570801765   0.9680547229935842   0.5938450129477865   0.6828163520584886   0.9129691528587722   0.7244865386403984   0.06232243195772163   0.27659311645494516   0.8104385526656283   0.16871870573393144   0.12451795438009036   0.12187405253673965   0.8726648930184753
0.4636909233459171   0.4454693126321418   0.6604074719397525   0.7502038445315969   0.4988768468130004   0.721239805320038   0.42645749224505286   0.5182059278228707   0.28570847643009356   0.6586092726266446   0.8750454208411573   0.08464197211485298   0.31765375343650937   0.06476425967885815   0.19222906878266868   0.17167281925608077   0.593167214796111   0.002441827721136534   0.9156359523277235   0.36123426659045255   0.4244485090621795   0.8779238733410462   0.7937618997909839   0.4885693735719772   0.9607575857162625   0.43245456070890437   0.13335442785123136   0.7383655290403802   0.46188073890326203   0.7112147553888665   0.7068969356061785   0.22015960121750958   0.1761722624731685   0.052605482762221795   0.8318515147650212   0.1355176291026566   0.8585185090366592   0.9878412230833636   0.6396224459823525   0.9638448098465758   0.26535129424054815   0.9853993953622271   0.7239864936546291   0.6026105432561233   0.8409027851783687   0.10747552202118094   0.9302245938636452   0.11404116968414608   0.8801451994621062   0.6750209613122765   0.7968701660124138   0.37567564064376585   0.4182644605588442   0.9638062059234102   0.08997323040623531   0.15551603942625628   0.24209219808567572   0.9112007231611883   0.2581217156412141   0.01999841032359967   0.38357368904901656   0.9233595000778246   0.6184992696588616   0.05615360047702385
0.11822239480846841   0.9379601047155975   0.8945127760042325   0.45354305722090055   0.2773196096300998   0.8304845826944166   0.9642881821405873   0.3395018875367545   0.39717441016799354   0.1554636213821401   0.1674180161281735   0.9638262468929886   0.9789099496091493   0.19165741545872997   0.07744478572193818   0.8083102074667323   0.7368177515234736   0.28045669229754167   0.8193230700807241   0.7883117971431327   0.353244062474457   0.357097192219717   0.20082380042186254   0.7321581966661088   0.2350216676659886   0.4191370875041194   0.30631102441763003   0.27861513944520827   0.9577020580358888   0.5886525048097028   0.3420228422770427   0.9391132519084538   0.5605276478678953   0.4331888834275626   0.1746048261488692   0.9752870050154652   0.581617698258746   0.24153146796883265   0.09716004042693102   0.16697679754873282   0.8447999467352724   0.961074775671291   0.2778369703462069   0.37866500040560014   0.49155588426081537   0.603977583451574   0.07701316992434441   0.6465068037394913   0.2565342165948268   0.18484049594745466   0.7707021455067143   0.367891664294283   0.29883215855893797   0.5961879911377519   0.4286793032296717   0.4287784123858292   0.7383045106910426   0.16299910771018927   0.2540744770808025   0.45349140737036403   0.15668681243229665   0.9214676397413566   0.15691443665387145   0.2865146098216312
0.3118868656970243   0.9603928640700656   0.8790774663076645   0.9078496094160311   0.8203309814362089   0.3564152806184916   0.8020642963833201   0.2613428056765398   0.5637967648413821   0.17157478467103693   0.031362150876605724   0.8934511413822568   0.2649646062824441   0.575386793533285   0.602682847646934   0.46467272899642753   0.5266600955914015   0.4123876858230957   0.34860837056613153   0.011181321626063504   0.3699732831591048   0.4909200460817391   0.1916939339122601   0.7246667118044323   0.058086417462080576   0.5305271820116735   0.3126164676045956   0.8168171023884012   0.2377554360258717   0.17411190139318192   0.5105521712212755   0.5554742967118614   0.6739586711844896   0.0025371167221449878   0.4791900203446698   0.6620231553296048   0.4089940649020455   0.42715032318886   0.8765071726977357   0.19735042633317718   0.882333969310644   0.014762637365764282   0.5278988021316041   0.18616910470711368   0.5123606861515392   0.5238425912840252   0.3362048682193441   0.46150239290268136   0.4542742686894585   0.9933154092723517   0.023588400614748484   0.6446852905142801   0.21651883266358685   0.8192035078791698   0.513036229393473   0.08921099380241868   0.5425601614790972   0.8166663911570248   0.03384620904880324   0.42718783847281394   0.1335660965770518   0.38951606796816485   0.15733903635106752   0.2298374121396368
0.2512321272664078   0.3747534306024005   0.6294402342194634   0.04366830743252312   0.7388714411148687   0.8509108393183753   0.2932353660001193   0.5821659145298418   0.28459717242541016   0.8575954300460237   0.2696469653853708   0.9374806240155616   0.0680783397618233   0.03839192216685383   0.7566107359918978   0.8482696302131429   0.5255181782827261   0.22172553100982903   0.7227645269430946   0.42108179174032895   0.39195208170567425   0.8322094630416642   0.5654254905920271   0.19124437960069215   0.14071995443926644   0.45745603243926364   0.9359852563725637   0.14757607216816904   0.40184851332439775   0.6065451931208883   0.6427498903724445   0.5654101576383272   0.11725134089898759   0.7489497630748646   0.3731029249870736   0.6279295336227657   0.0491730011371643   0.7105578409080108   0.6164921889951759   0.7796599034096228   0.5236548228544382   0.4888323098981818   0.8937276620520813   0.3585781116692938   0.13170274114876399   0.6566228468565176   0.32830217146005425   0.16733373206860166   0.9909827867094976   0.19916681441725395   0.39231691508749056   0.019757659900432607   0.5891342733850998   0.5926216212963656   0.7495670247150462   0.4543475022621053   0.47188293248611224   0.843671858221501   0.37646409972797257   0.8264179686393396   0.4227099313489479   0.1331140173134902   0.7599719107327967   0.04675806522971682
0.8990551084945096   0.6442817074153084   0.8662442486807155   0.688179953560423   0.7673523673457456   0.9876588605587908   0.5379420772206612   0.5208462214918214   0.7763695806362481   0.7884920461415368   0.1456251621331706   0.5010885615913887   0.1872353072511483   0.19587042484517114   0.39605813741812446   0.04674105932928343   0.7153523747650361   0.35219856662367016   0.019594037690151882   0.22032309068994382   0.29264244341608814   0.21908454931017993   0.25962212695735515   0.173565025460227   0.39358733492157844   0.5748028418948715   0.3933778782766397   0.485385071899804   0.6262349675758327   0.5871439813360808   0.8554358010559786   0.9645388504079827   0.8498653869395847   0.7986519351945439   0.7098106389228079   0.46345028881659395   0.6626300796884363   0.6027815103493728   0.31375250150468353   0.4167092294873105   0.9472777049234004   0.25058294372570267   0.29415846381453165   0.1963861387973667   0.6546352615073122   0.03149839441552272   0.034536336857176476   0.022821113337139678   0.2610479265857337   0.4566955525206512   0.6411584585805368   0.5374360414373357   0.634812959009901   0.8695515711845704   0.7857226575245582   0.572897191029353   0.7849475720703163   0.07089963599002647   0.07591201860175023   0.10944690221275907   0.12231749238187987   0.4681181256406537   0.7621595170970668   0.6927376727254486
0.17503978745847953   0.21753518191495103   0.46800105328253505   0.4963515339280819   0.5204045259511674   0.1860367874994283   0.4334647164253586   0.4735304205909422   0.25935659936543365   0.7293412349787771   0.7923062578448219   0.9360943791536065   0.6245436403555327   0.8597896637942067   0.006583600320263664   0.36319718812425356   0.8395960682852164   0.7888900278041803   0.9306715817185134   0.25375028591149446   0.7172785759033365   0.3207719021635266   0.16851206462144672   0.5610126131860459   0.542238788444857   0.10323672024857555   0.7005110113389117   0.06466107925796402   0.021834262493689652   0.9171999327491472   0.26704629491355303   0.5911306586670219   0.762477663128256   0.18785869777037012   0.4747400370687312   0.6550362795134153   0.13793402277272335   0.3280690339761634   0.4681564367484675   0.29183909138916175   0.29833795448750694   0.5391790061719831   0.5374848550299541   0.03808880547766729   0.5810593785841703   0.21840710400845656   0.3689727904085074   0.4770761922916214   0.03882059013931337   0.11517038375988102   0.6684617790695957   0.41241511303365735   0.016986327645623717   0.19797045101073377   0.40141548415604267   0.8212844543666356   0.2545086645173677   0.010111753240363655   0.9266754470873115   0.16624817485322027   0.11657464174464434   0.6820427192642002   0.45851901033884396   0.8744090834640585
0.8182366872571374   0.14286371309221713   0.9210341553088899   0.8363202779863912   0.23717730867296705   0.9244566090837606   0.5520613649003825   0.35924408569476984   0.19835671853365366   0.8092862253238795   0.8835995858307867   0.9468289726611124   0.18137039088802998   0.6113157743131458   0.482184101674744   0.12554451829447688   0.9268617263706622   0.6012040210727821   0.5555086545874326   0.9592963434412566   0.810287084626018   0.9191613018085818   0.0969896442485886   0.08488725997719809   0.9920503973688806   0.7762975887163647   0.17595548893969876   0.24856698199080687   0.7548730886959135   0.8518409796326042   0.6238941240393163   0.889322896296037   0.5565163701622597   0.04255475430872466   0.7402945382085295   0.9424939236349246   0.3751459792742298   0.4312389799955789   0.2581104365337855   0.8169494053404477   0.44828425290356755   0.8300349589227968   0.7026017819463529   0.8576530618991911   0.6379971682775496   0.910873657114215   0.6056121376977643   0.772765801921993   0.6459467709086691   0.13457606839785025   0.4296566487580656   0.5241988199311861   0.8910736822127556   0.28273508876524606   0.8057625247187493   0.6348759236351491   0.3345573120504958   0.2401803344565214   0.06546798651021977   0.6923820000002245   0.959411332776266   0.8089413544609425   0.8073575499764343   0.8754325946597769
0.5111270798726985   0.9789063955381457   0.1047557680300813   0.017779532760585783   0.8731299115951489   0.0680327384239307   0.49914363033231696   0.24501373083859282   0.22718314068647974   0.9334566700260805   0.06948698157425133   0.7208149109074067   0.3361094584737241   0.6507215812608343   0.263724456855502   0.08593898727225763   0.0015521464232282531   0.410541246804313   0.19825647034528224   0.3935569872720331   0.04214081364696224   0.6015998923433705   0.390898920368848   0.5181243926122563   0.5310137337742638   0.6226934968052248   0.2861431523387667   0.5003448598516705   0.6578838221791149   0.554660758381294   0.7869995220064497   0.2553311290130777   0.43070068149263524   0.6212040883552137   0.7175125404321984   0.534516218105671   0.09459122301891112   0.9704825070943792   0.4537880835766964   0.44857723083341333   0.09303907659568288   0.5599412602900663   0.25553161323141416   0.05502024356138024   0.05089826294872063   0.9583413679466958   0.8646326928625662   0.536895850949124   0.5198845291744568   0.335647871141471   0.5784895405237995   0.036550991097453474   0.8620007069953419   0.780987112760177   0.7914900185173498   0.7812198620843758   0.4313000255027067   0.15978302440496328   0.07397747808515137   0.24670364397870484   0.33670880248379553   0.18930051731058406   0.620189394508455   0.7981264131452915
0.24366972588811267   0.6293592570205178   0.3646577812770408   0.7431061695839113   0.19277146293939204   0.671017889073822   0.5000250884144746   0.20621031863478728   0.6728869337649352   0.335370017932351   0.9215355478906752   0.16965932753733381   0.8108862267695933   0.5543829051721741   0.13004552937332534   0.388439465452958   0.37958620126688664   0.3945998807672108   0.05606805128817397   0.14173582147425318   0.04287739878309108   0.20529936345662678   0.435878656779719   0.3436094083289617   0.7992076728949784   0.5759401064361089   0.07122087550267821   0.6005032387450504   0.6064362099555863   0.904922217362287   0.5711957870882036   0.3942929201102631   0.9335492761906512   0.569552199429936   0.6496602391975285   0.22463359257292934   0.12266304942105787   0.01516929425776185   0.5196147098242031   0.8361941271199713   0.7430768481541712   0.6205694134905511   0.46354665853602917   0.6944583056457181   0.7001994493710801   0.41527005003392425   0.027668001756310175   0.35084889731675645   0.9009917764761017   0.8393299435978153   0.9564471262536319   0.750345658571706   0.29455556652051534   0.9344077262355284   0.38525133916542836   0.35605273846144286   0.3610062903298642   0.36485552680559236   0.7355910999678998   0.13141914588851356   0.23834324090880635   0.3496862325478305   0.21597639014369674   0.29522501876854224
0.49526639275463513   0.7291168190572794   0.7524297316076676   0.600766713122824   0.795066943383555   0.31384676902335523   0.7247617298513573   0.24991781580606764   0.8940751669074533   0.4745168254255399   0.7683146035977254   0.4995721572343616   0.5995196003869379   0.5401090991900116   0.38306326443229705   0.14351941877291874   0.23851331005707366   0.17525357238441924   0.6474721644643971   0.012100272884405194   0.00017006914826731088   0.8255673398365887   0.4314957743207004   0.716875254115863   0.5049036763936322   0.09645052077930925   0.6790660427130328   0.11610854099303887   0.7098367330100772   0.7826037517559541   0.9543043128616754   0.8661907251869713   0.8157615661026241   0.3080869263304141   0.18598970926395003   0.3666185679526096   0.21624196571568619   0.7679778271404025   0.802926444831653   0.22309914917969087   0.9777286556586126   0.5927242547559832   0.15545428036725584   0.2109988762952857   0.9775585865103452   0.7671569149193945   0.7239585060465554   0.49412362217942274   0.472654910116713   0.6707063941400853   0.044892463333522606   0.37801508118638383   0.7628181771066358   0.8881026423841312   0.09058815047184716   0.5118243559994126   0.9470566110040117   0.580015716053717   0.9045984412078971   0.14520578804680298   0.7308146452883255   0.8120378889133146   0.10167199637624418   0.9221066388671121
0.7530859896297131   0.21931363415733132   0.9462177160089883   0.7111077625718264   0.7755274031193679   0.4521567192379368   0.2222592099624329   0.2169841403924037   0.30287249300265484   0.7814503250978515   0.17736674662891028   0.8389690592060198   0.540054315896019   0.8933476827137203   0.08677859615706311   0.32714470320660727   0.5929977048920073   0.31333196666000324   0.18218015494916595   0.18193891515980426   0.8621830596036818   0.5012940777466887   0.08050815857292179   0.2598322762926922   0.10909706997396872   0.2819804435893573   0.13429044256393347   0.5487245137208657   0.3335696668546009   0.8298237243514205   0.9120312326015005   0.331740373328462   0.03069717385194606   0.048373399253569   0.7346644859725903   0.4927713141224422   0.490642857955927   0.15502571653984867   0.6478858898155272   0.16562661091583492   0.8976451530639197   0.8416937498798455   0.4657057348663612   0.9836876957560307   0.035462093460237924   0.3403996721331568   0.3851975762934394   0.7238554194633385   0.9263650234862693   0.058419228543799495   0.25090713372950596   0.17513090574247275   0.5927953566316684   0.22859550419237898   0.33887590112800536   0.8433905324140107   0.5620981827797222   0.18022210493880997   0.6042114151554151   0.35061921829156856   0.07145532482379527   0.0251963883989613   0.9563255253398879   0.18499260737573367
0.1738101717598756   0.18350263851911586   0.4906197904735267   0.20130491161970301   0.13834807829963766   0.843102966385959   0.10542221418008732   0.4774494921563645   0.21198305481336846   0.7846837378421595   0.8545150804505813   0.30231858641389175   0.6191876981817002   0.5560882336497806   0.515639179322576   0.458928053999881   0.05708951540197787   0.3758661287109706   0.9114277641671609   0.10830883570831246   0.9856341905781826   0.35066974031200926   0.955102238827273   0.9233162283325788   0.811824018818307   0.16716710179289343   0.4644824483537462   0.7220113167128758   0.6734759405186693   0.3240641354069344   0.3590602341736589   0.24456182455651124   0.4614928857053009   0.5393803975647748   0.5045451537230775   0.9422432381426195   0.8423051875236007   0.9832921639149943   0.9889059744005015   0.48331518414273844   0.7852156721216229   0.6074260352040237   0.07747821023334069   0.375006348434426   0.7995814815434403   0.25675629489201446   0.12237597140606775   0.45169012010184717   0.9877574627251333   0.08958919309912101   0.6578935230523215   0.7296788033889714   0.31428152220646394   0.7655250576921866   0.2988332888786626   0.48511697883246013   0.852788636501163   0.22614466012741175   0.7942881351555852   0.5428737406898407   0.01048344897756227   0.24285249621241742   0.8053821607550835   0.05955855654710227
0.22526777685593938   0.6354264610083937   0.7279039505217428   0.6845522081126764   0.4256862953124991   0.37867016611637927   0.6055279791156751   0.23286208801082914   0.4379288325873658   0.2890809730172582   0.9476344560633536   0.5031832846218578   0.12364731038090186   0.5235559153250716   0.6488011671846909   0.0180663057893976   0.27085867387973883   0.2974112551976599   0.8545130320291059   0.47519256509955693   0.26037522490217657   0.054558758985242456   0.049130871274022284   0.41563400855245464   0.035107448046237194   0.41913229797684876   0.32122692075227943   0.7310818004397783   0.6094211527337381   0.04046213186046952   0.7156989416366043   0.4982197124289492   0.1714923201463723   0.7513811588432113   0.7680644855732507   0.9950364278070915   0.047845009765470445   0.22782524351813968   0.11926331838855975   0.9769701220176938   0.7769863358857316   0.9304139883204798   0.2647502863594539   0.5017775569181369   0.516611110983555   0.8758552293352373   0.21561941508543164   0.08614354836568228   0.48150366293731783   0.4567229313583886   0.8943924943331523   0.35506174792590395   0.8720825102035797   0.41626079949791905   0.17869355269654794   0.8568420354969548   0.7005901900572075   0.6648796406547077   0.4106290671232972   0.8618056076898634   0.652745180291737   0.4370543971365681   0.2913657487347375   0.8848354856721695
0.8757588444060054   0.5066404088160883   0.026615462375283564   0.3830579287540326   0.3591477334224503   0.630785179480851   0.810996047289852   0.29691438038835033   0.8776440704851325   0.1740622481224624   0.9166035529566997   0.9418526324624464   0.005561560281552717   0.7578014486245434   0.7379100002601517   0.08501059696549162   0.3049713702243453   0.09292180796983558   0.3272809331368545   0.2232049892756283   0.6522261899326083   0.6558674108332675   0.03591518440211706   0.33836950360345874   0.7764673455266029   0.14922700201717917   0.009299722026833499   0.9553115748494262   0.41731961210415264   0.5184418225363282   0.19830367473698157   0.6583971944610758   0.5396755416190202   0.3443795744138658   0.28170012178028186   0.7165445619986294   0.5341139813374675   0.5865781257893224   0.5437901215201301   0.6315339650331377   0.22914261111312217   0.4936563178194869   0.21650918838327554   0.4083289757575095   0.5769164211805139   0.8377889069862194   0.1805940039811585   0.06995947215405074   0.8004490756539109   0.6885619049690402   0.171294281954325   0.1146478973046246   0.38312946354975824   0.170120082432712   0.9729906072173434   0.4562507028435488   0.8434539219307381   0.8257405080188462   0.6912904854370615   0.7397061408449194   0.30933994059327063   0.2391623822295237   0.14750036391693147   0.1081721758117816
0.08019732948014847   0.7455060644100368   0.930991175533656   0.6998432000542721   0.5032809082996347   0.9077171574238174   0.7503971715524974   0.6298837279002213   0.7028318326457237   0.21915525245477716   0.5791028895981725   0.5152358305955967   0.31970236909596544   0.04903517002206514   0.606112282380829   0.058985127752047964   0.47624844716522735   0.22329466200321896   0.9148217969437674   0.3192789869071286   0.16690850657195672   0.9841322797736952   0.767321433026836   0.21110681109534699   0.08671117709180824   0.23862621536365844   0.8363302574931801   0.5112636110410749   0.5834302687921736   0.33090905793984104   0.08593308594068265   0.8813798831408536   0.88059843614645   0.11175380548506389   0.5068301963425103   0.36614405254525684   0.5608960670504844   0.06271863546299876   0.9007179139616812   0.30715892479320883   0.08464761988525708   0.8394239734597798   0.9858961170179137   0.9878799378860803   0.9177391133133004   0.8552916936860846   0.2185746839910777   0.7767731267907333   0.8310279362214921   0.6166654783224261   0.38224442649789764   0.26550951574965836   0.2475976674293185   0.2857564203825851   0.296311340557215   0.3841296326088048   0.3669992312828686   0.1740026148975212   0.7894811442147048   0.017985580063547987   0.8061031642323842   0.11128397943452244   0.8887632302530236   0.7108266552703392
0.7214555443471271   0.27186000597474264   0.9028671132351099   0.7229467173842589   0.8037164310338267   0.41656831228865804   0.6842924292440322   0.9461735905935256   0.9726884948123347   0.799902833966232   0.3020480027461345   0.6806640748438673   0.7250908273830161   0.5141464135836469   0.005736662188919538   0.2965344422350624   0.3580915961001475   0.34014379868612565   0.21625551797421474   0.2785488621715144   0.5519884318677634   0.22885981925160323   0.32749228772119116   0.5677222069011753   0.8305328875206364   0.9569998132768606   0.4246251744860812   0.8447754895169164   0.02681645648680961   0.5404315009882026   0.7403327452420491   0.8986018989233908   0.054127961674475006   0.7405286670219706   0.43828474249591454   0.2179378240795236   0.32903713429145887   0.22638225343832374   0.432548080306995   0.9214033818444612   0.9709455381913114   0.8862384547521981   0.21629256233278027   0.6428545196729467   0.418957106323548   0.6573786355005948   0.8888002746115892   0.07513231277177146   0.5884242188029116   0.7003788222237343   0.4641751001255079   0.23035682325485501   0.561607762316102   0.15994732123553168   0.7238423548834588   0.33175492433146414   0.507479800641627   0.41941865421356106   0.28555761238754424   0.11381710025194054   0.17844266635016814   0.19303640077523732   0.8530095320805492   0.19241371840747934
0.2074971281588568   0.3067979460230392   0.6367169697477689   0.5495591987345326   0.7885400218353088   0.6494193105224444   0.7479166951361799   0.4744268859627611   0.20011580303239718   0.9490404882987101   0.283741595010672   0.24407006270790613   0.6385080407162952   0.7890931670631784   0.5598992401272131   0.912315138376442   0.13102824007466812   0.3696745128496174   0.27434162773966897   0.7984980381245014   0.9525855737244999   0.17663811207438004   0.4213320956591197   0.606084319717022   0.7450884455656431   0.8698401660513408   0.7846151259113507   0.05652512098248948   0.9565484237303343   0.22042085552889643   0.036698430775170876   0.5820982350197283   0.7564326206979372   0.27138036723018627   0.7529568357644989   0.33802817231182225   0.11792457998164202   0.4822872001670078   0.1930575956372857   0.4257130339353803   0.9868963399069739   0.11261268731739045   0.9187159678976168   0.6272149958108789   0.03431076618247394   0.9359745752430104   0.497383872238497   0.02113067609385681   0.2892223206168308   0.06613440919166957   0.7127687463271463   0.9646055551113674   0.3326738968864964   0.8457135536627731   0.6760703155519754   0.382507320091639   0.5762412761885592   0.5743331864325868   0.9231134797874765   0.04447914777981676   0.45831669620691723   0.09204598626557901   0.7300558841501908   0.6187661138444365
0.47142035629994333   0.9794332989481885   0.8113399162525741   0.9915511180335577   0.4371095901174694   0.04345872370517817   0.31395604401407706   0.9704204419397008   0.14788726950063863   0.9773243145135087   0.6011872976869308   0.005814886828333477   0.8152133726141422   0.13161076085073545   0.9251169821349554   0.6233075667366945   0.23897209642558295   0.5572775744181486   0.002003502347478838   0.5788284189568778   0.7806554002186658   0.4652315881525696   0.271947618197288   0.9600623051124413   0.30923504391872236   0.485798289204381   0.4606077019447139   0.9685111870788836   0.872125453801253   0.44233956549920284   0.1466516579306368   0.9980907451391828   0.7242381843006143   0.46501525098569424   0.545464360243706   0.9922758583108493   0.9090248116864721   0.3334044901349588   0.6203473781087506   0.36896829157415484   0.6700527152608892   0.7761269157168101   0.6183438757612718   0.7901398726172771   0.8893973150422234   0.3108953275642406   0.34639625756398384   0.8300775675048359   0.580162271123501   0.8250970383598596   0.88578855561927   0.8615663804259522   0.7080368173222481   0.3827574728606567   0.7391368976886331   0.8634756352867695   0.9837986330216338   0.9177422218749625   0.19367253744492707   0.8711997769759201   0.07477382133516174   0.5843377317400037   0.5733251593361764   0.5022314854017653
0.4047211060742726   0.8082108160231934   0.9549812835749045   0.7120916127844882   0.5153237910320492   0.4973154884589529   0.6085850260109208   0.8820140452796523   0.935161519908548   0.6722184500990933   0.7227964703916508   0.020447664853700035   0.2271247025862999   0.28946097723843656   0.9836595727030177   0.15697202956693057   0.24332606956466607   0.3717187553634741   0.7899870352580907   0.2857722525910104   0.16855224822950435   0.7873810236234704   0.21666187592191422   0.7835407671892451   0.7638311421552317   0.979170207600277   0.26168059234700963   0.07144915440475694   0.24850735112318262   0.48185471914132405   0.6530955663360889   0.18943510912510464   0.3133458312146346   0.8096362690422307   0.930299095944438   0.1689874442714046   0.08622112862833468   0.5201752918037942   0.9466395232414204   0.012015414704474035   0.8428950590636686   0.14845653644032009   0.15665248798332979   0.7262431621134636   0.6743428108341643   0.36107551281684963   0.9399906120614155   0.9427023949242185   0.9105116686789325   0.3819053052165727   0.678310019714406   0.8712532405194615   0.6620043175557498   0.9000505860752486   0.025214453378317046   0.6818181313943569   0.3486584863411153   0.09041431703301785   0.09491535743387897   0.5128306871229523   0.2624373577127806   0.5702390252292237   0.14827583419245857   0.5008152724184782
0.419542298649112   0.42178248878890356   0.9916233462091287   0.7745721103050146   0.7451994878149477   0.06070697597205391   0.05163273414771321   0.8318697153807961   0.8346878191360152   0.6788016707554813   0.3733227144333073   0.9606164748613346   0.17268350158026535   0.7787510846802326   0.3481082610549902   0.27879834346697774   0.8240250152391501   0.6883367676472147   0.25319290362111124   0.7659676563440254   0.5615876575263694   0.11809774241799112   0.1049170694286527   0.26515238392554713   0.14204535887725742   0.6963152536290875   0.11329372321952391   0.49058027362053247   0.3968458710623097   0.6356082776570336   0.06166098907181071   0.6587105582397363   0.5621580519262944   0.9568066069015524   0.6883382746385034   0.6980940833784017   0.3894745503460291   0.17805552222131982   0.34023001358351324   0.41929573991142394   0.5654495351068791   0.4897187545741051   0.08703710996240195   0.6533280835673986   0.00386187758050964   0.37162101215611393   0.9821200405337492   0.3881756996418514   0.8618165187032523   0.6753057585270263   0.8688263173142253   0.8975954260213189   0.46497064764094254   0.03969748086999275   0.8071653282424146   0.23888486778158258   0.9028125957146481   0.08289087396844033   0.11882705360391119   0.5407907844031808   0.5133380453686189   0.9048353517471205   0.778597040020398   0.12149504449175692
0.9478885102617399   0.41511659717301547   0.691559930057996   0.4681669609243584   0.9440266326812302   0.04349558501690151   0.7094398895242467   0.079991261282507   0.08221011397797803   0.36818982648987514   0.8406135722100214   0.1823958352611881   0.6172394663370355   0.3284923456198824   0.03344824396760683   0.9435109674796055   0.7144268706223874   0.24560147165144205   0.9146211903636956   0.40272018307642465   0.20108882525376845   0.34076611990432154   0.13602415034329768   0.28122513858466774   0.25320031499202855   0.9256495227313061   0.44446422028530164   0.8130581776603093   0.3091736823107983   0.8821539377144045   0.7350243307610549   0.7330669163778023   0.22696356833282028   0.5139641112245295   0.8944107585510335   0.5506710811166142   0.6097241019957848   0.18547176560464707   0.8609625145834265   0.6071601136370087   0.8952972313733973   0.939870293953205   0.9463413242197309   0.20443993056058404   0.6942084061196289   0.5991041740488835   0.8103171738764333   0.9232147919759163   0.4410080911276003   0.6734546513175774   0.3658529535911316   0.110156614315607   0.131834408816802   0.7913007136031729   0.6308286228300768   0.37708969793780467   0.9048708404839817   0.2773366023786434   0.7364178642790433   0.8264186168211904   0.295146738488197   0.09186483677399632   0.8754553496956168   0.21925850318418177
0.39984950711479966   0.15199454282079128   0.9291140254758858   0.014818572623597722   0.7056411009951707   0.5528903687719078   0.11879685159945254   0.0916037806476814   0.2646330098675705   0.8794357174543304   0.752943898008321   0.9814471663320744   0.13279860105076846   0.08813500385115754   0.12211527517824415   0.6043574683942697   0.2279277605667867   0.8107984014725141   0.38569741089920084   0.7779388515730793   0.9327810220785897   0.7189335646985179   0.5102420612035841   0.5586803483888976   0.5329315149637901   0.5669390218777266   0.5811280357276982   0.5438617757652998   0.8272904139686192   0.014048653105818765   0.46233118412824575   0.4522579951176184   0.5626574041010488   0.13461293565148838   0.7093872861199249   0.470810828785544   0.42985880305028035   0.04647793180033084   0.5872720109416807   0.8664533603912743   0.20193104248349364   0.2356795303278167   0.20157460004247985   0.08851450881819498   0.26915002040490393   0.5167459656292989   0.6913325388388958   0.5298341604292974   0.7362185054411139   0.9498069437515723   0.11020450311119752   0.9859723846639976   0.9089280914724946   0.9357582906457536   0.6478733189829518   0.5337143895463793   0.34627068737144584   0.8011453549942652   0.9384860328630269   0.06290356076083525   0.9164118843211655   0.7546674231939343   0.35121402192134626   0.19645020036956098
0.7144808418376718   0.5189878928661176   0.14963942187886642   0.10793569155136601   0.4453308214327679   0.002241927236818755   0.45830688303997064   0.5781015311220685   0.709112315991654   0.05243498348524645   0.34810237992877313   0.5921291464580709   0.8001842245191594   0.11667669283949292   0.7002290609458214   0.058414756911691665   0.4539135371477136   0.31553133784522774   0.7617430280827944   0.9955111961508564   0.5375016528265482   0.5608639146512935   0.4105290061614481   0.7990609957812954   0.8230208109888763   0.04187602178517583   0.2608895842825817   0.6911253042299295   0.37768998955610833   0.039634094548357084   0.802582701242611   0.11302377310786084   0.6685776735644543   0.9871991110631106   0.4544803213138379   0.5208946266497899   0.8683934490452949   0.8705224182236178   0.7542512603680166   0.4624798697380983   0.41447991189758127   0.55499108037839   0.9925082322852222   0.46696867358724187   0.8769782590710331   0.9941271657270965   0.5819792261237741   0.6679076778059464   0.05395744808215684   0.9522511439419207   0.32108964184119243   0.976782373576017   0.6762674585260485   0.9126170493935636   0.5185069405985814   0.8637586004681562   0.007689784961594179   0.9254179383304529   0.06402661928474344   0.34286397381836625   0.1392963359162993   0.054895520106835245   0.30977535891672686   0.880384104080268
0.724816424018718   0.4999044397284453   0.31726712663150464   0.4134154304930261   0.8478381649476849   0.5057772740013488   0.7352879005077305   0.7455077526870797   0.7938807168655281   0.5535261300594281   0.41419825866653814   0.7687253791110626   0.11761325833947961   0.6409090806658645   0.8956913180679568   0.9049667786429064   0.10992347337788543   0.7154911423354116   0.8316646987832134   0.5621028048245402   0.9706271374615861   0.6605956222285763   0.5218893398664864   0.6817187007442722   0.24581071344286806   0.160691182500131   0.20462221323498184   0.2683032702512461   0.39797254849518315   0.6549139084987823   0.4693343127272513   0.5227955175641664   0.6040918316296551   0.10138777843935415   0.05513605406071316   0.7540701384531038   0.4864785732901754   0.46047869777348965   0.1594447359927564   0.8491033598101974   0.37655509991228997   0.744987555438078   0.3277800372095431   0.28700055498565713   0.4059279624507039   0.0843919332095018   0.8058906973430566   0.6052818542413849   0.1601172490078358   0.9237007507093707   0.6012684841080748   0.3369785839901388   0.7621447005126527   0.2687868422105885   0.13193417138082347   0.8141830664259724   0.15805286888299766   0.16739906377123437   0.07679811732011031   0.06011292797286857   0.6715742955928222   0.7069203659977448   0.9173533813273539   0.21100956816267125
0.29501919568053225   0.9619328105596666   0.5895733441178108   0.9240090131770141   0.8890912332298283   0.8775408773501648   0.7836826467747542   0.31872715893562925   0.7289739842219926   0.9538401266407941   0.18241416266667948   0.9817485749454905   0.9668292837093398   0.6850532844302055   0.050479991285856   0.1675655085195181   0.8087764148263422   0.5176542206589712   0.9736818739657457   0.10745258054664954   0.13720211923351996   0.8107338546612265   0.05632849263839177   0.8964430123839783   0.8421829235529877   0.8488010441015598   0.4667551485205809   0.9724339992069642   0.9530916903231594   0.9712601667513949   0.6830725017458267   0.653706840271335   0.22411770610116685   0.017420040110600887   0.5006583390791473   0.6719582653258445   0.25728842239182703   0.33236675568039536   0.4501783477932912   0.5043927568063263   0.4485120075654848   0.8147125350214242   0.4764964738275455   0.39694017625967687   0.3113098883319648   0.0039786803601977215   0.42016798118915377   0.5004971638756985   0.4691269647789771   0.15517763625863792   0.9534128326685728   0.5280631646687344   0.5160352744558176   0.18391746950724297   0.2703403309227461   0.8743563243973994   0.2919175683546508   0.16649742939664208   0.769681991843599   0.20239805907155495   0.03462914596282382   0.8341306737162467   0.31950364405030773   0.6980053022652285
0.586117138397339   0.01941813869482257   0.8430071702227622   0.3010651260055517   0.27480725006537415   0.015439458334624848   0.42283918903360845   0.8005679621298532   0.8056802852863971   0.8602618220759869   0.4694263563650356   0.2725047974611188   0.28964501083057936   0.6763443525687439   0.19908602544228948   0.3981484730637193   0.9977274424759286   0.5098469231721019   0.42940403359869056   0.1957504139921644   0.9630982965131047   0.6757162494558552   0.10990038954838283   0.49774511172693586   0.3769811581157657   0.6562981107610326   0.26689321932562066   0.19667998572138415   0.10217390805039155   0.6408586524264077   0.8440540302920122   0.39611202359153097   0.2964936227639945   0.7805968303504208   0.37462767392697655   0.12360722613041222   0.006848611933415076   0.10425247778167684   0.17554164848468706   0.7254587530666929   0.009121169457486521   0.5944055546095749   0.7461376148859965   0.5297083390745285   0.04602287294438179   0.9186893051537198   0.6362372253376136   0.031963227347592674   0.6690417148286161   0.26239119439268715   0.369344006011993   0.8352832416262085   0.5668678067782246   0.6215325419662794   0.5252899757199808   0.43917121803467757   0.2703741840142301   0.8409357116158586   0.15066230179300433   0.3155639919042653   0.26352557208081495   0.7366832338341818   0.9751206533083172   0.5901052388375724
0.2544044026233285   0.14227767922460682   0.22898303842232073   0.06039689976304391   0.20838152967894666   0.22358837407088705   0.5927458130847071   0.02843367241545124   0.5393398148503306   0.9611971796781998   0.223401807072714   0.1931504307892427   0.9724720080721061   0.33966463771192046   0.6981118313527331   0.7539792127545651   0.702097824057876   0.49872892609606184   0.5474495295597288   0.4384152208502998   0.43857225197706107   0.7620456922618801   0.5723288762514116   0.8483099820127274   0.1841678493537326   0.6197680130372732   0.34334583782909084   0.7879130822496835   0.9757863196747859   0.3961796389663862   0.7506000247443838   0.7594794098342322   0.43644650482445535   0.43498245928818635   0.5271982176716697   0.5663289790449896   0.46397449675234925   0.09531782157626591   0.8290863863189366   0.8123497662904244   0.7618766726944732   0.5965888954802041   0.28163685675920774   0.37393454544012455   0.32330442071741217   0.834543203218324   0.7093079805077962   0.5256245634273972   0.13913657136367957   0.21477519018105073   0.36596214267870536   0.7377114811777137   0.16335025168889364   0.8185955512146645   0.6153621179343216   0.9782320713434813   0.7269037468644383   0.38361309192647813   0.08816390026265182   0.41190309229849176   0.26292925011208906   0.28829527035021224   0.25907751394371525   0.5995533260080673
0.5010525774176159   0.6917063748700082   0.9774406571845075   0.2256187805679428   0.17774815670020372   0.8571631716516842   0.2681326766767113   0.6999942171405457   0.03861158533652414   0.6423879814706335   0.902170533998006   0.962282735962832   0.8752613336476305   0.8237924302559689   0.2868084160636844   0.9840506646193506   0.1483575867831922   0.4401793383294908   0.19864451580103257   0.5721475723208589   0.8854283366711031   0.15188406797927856   0.9395670018573173   0.9725942463127916   0.38437575925348727   0.46017769310927037   0.9621263446728099   0.7469754657448487   0.20662760255328355   0.6030145214575862   0.6939936679960985   0.04698124860430306   0.1680160172167594   0.9606265399869527   0.7918231339980926   0.08469851264147103   0.2927546835691289   0.13683410973098378   0.5050147179344082   0.10064784802212036   0.1443970967859367   0.696654771401493   0.3063702021333756   0.5285002757012615   0.2589687601148336   0.5447707034222145   0.3668032002760583   0.5559060293884699   0.8745930008613464   0.08459301031294403   0.40467685560324845   0.8089305636436213   0.6679653983080628   0.4815784888553578   0.7106831876071499   0.7619493150393182   0.4999493810913034   0.5209519488684051   0.9188600536090573   0.6772508023978471   0.2071946975221745   0.3841178391374213   0.4138453356746491   0.5766029543757267
0.06279760073623779   0.6874630677359284   0.10747513354127344   0.0481026786744653   0.8038288406214043   0.1426923643137139   0.7406719332652152   0.4921966492859954   0.9292358397600579   0.05809935400076989   0.3359950776619667   0.6832660856423741   0.261270441451995   0.5765208651454121   0.6253118900548168   0.9213167706030561   0.7613210603606917   0.05556891627700699   0.7064518364457595   0.24406596820520893   0.5541263628385171   0.6714510771395857   0.29260650077111044   0.6674630138294821   0.4913287621022793   0.9839880094036574   0.185131367229837   0.6193603351550169   0.6874999214808751   0.8412956450899435   0.44445943396462184   0.1271636858690215   0.7582640817208173   0.7831962910891735   0.10846435630265515   0.4438976002266473   0.49699364026882226   0.20667542594376148   0.4831524662478383   0.5225808296235913   0.7356725799081306   0.1511065096667545   0.7767006298020788   0.2785148614183824   0.18154621706961346   0.4796554325271688   0.4840941290309684   0.6110518475889002   0.6902174549673341   0.4956674231235114   0.29896276180113135   0.9916915124338833   0.002717533486458986   0.6543717780335679   0.8545033278365095   0.8645278265648618   0.24445345176564168   0.8711754869443944   0.7460389715338543   0.42063022633821456   0.7474598114968194   0.664500061000633   0.26288650528601604   0.8980493967146232
0.011787231588688822   0.5133935513338784   0.4861858754839372   0.6195345352962409   0.8302410145190754   0.033738118806709606   0.002091746452968877   0.008482687707340675   0.14002355955174123   0.5380706956831982   0.7031289846518375   0.016791175273457325   0.13730602606528222   0.8836989176496302   0.848625656815328   0.15226334870859545   0.8928525742996405   0.012523430705235773   0.10258668528147363   0.7316331223703809   0.1453927628028211   0.34802336970460285   0.8397001799954575   0.8335837256557577   0.13360553121413227   0.8346298183707245   0.3535143045115204   0.21404919035951678   0.30336451669505693   0.8008916995640148   0.3514225580585515   0.2055665026521761   0.16334095714331573   0.26282100388081664   0.648293573406714   0.18877532737871877   0.02603493107803349   0.3791220862311865   0.7996679165913859   0.03651197867012331   0.13318235677839296   0.3665986555259507   0.6970812313099123   0.3048788562997424   0.9877895939755719   0.01857528582134785   0.8573810513144547   0.47129513064398476   0.8541840627614395   0.1839454674506234   0.5038667468029344   0.25724594028446796   0.5508195460663826   0.38305376788660855   0.1524441887443829   0.05167943763229189   0.3874785889230669   0.12023276400579191   0.5041506153376689   0.8629041102535732   0.3614436578450334   0.7411106777746055   0.704482698746283   0.8263921315834498
0.22826130106664047   0.3745120222486547   0.00740146743637063   0.5215132752837074   0.24047170709106863   0.3559367364273069   0.15002041612191588   0.05021814463972267   0.38628764432962903   0.17199126897668346   0.6461536693189815   0.7929722043552547   0.8354680982632464   0.7889375010900749   0.4937094805745986   0.7412927667229628   0.4479895093401795   0.668704737084283   0.9895588652369297   0.8783886564693897   0.08654585149514607   0.9275940593096775   0.2850761664906467   0.05199652488593987   0.8582845504285056   0.5530820370610228   0.27767469905427605   0.5304832496022325   0.617812843337437   0.19714530063371594   0.12765428293236017   0.4802651049625098   0.2315251990078079   0.025154031657032484   0.4815006136133787   0.6872929006072551   0.3960571007445615   0.2362165305669576   0.9877911330387801   0.9460001338842923   0.948067591404382   0.5675117934826747   0.9982322678018504   0.06761147741490262   0.861521739909236   0.6399177341729971   0.7131561013112037   0.01561495252896274   0.0032371894807303268   0.08683569711197427   0.43548140225692766   0.4851317029267303   0.38542434614329335   0.8896903964782583   0.30782711932456747   0.004866597964220487   0.15389914713548544   0.8645363648212259   0.8263265057111888   0.3175736973569654   0.7578420463909239   0.6283198342542682   0.8385353726724087   0.37157356347267306
0.8097744549865419   0.06080804077159361   0.8403031048705583   0.3039620860577705   0.948252715077306   0.42089030659859655   0.12714700355935457   0.28834713352880775   0.9450155255965756   0.33405460948662224   0.6916656013024269   0.8032154306020775   0.5595911794532823   0.44436421300836393   0.38383848197785947   0.7983488326378569   0.4056920323177969   0.5798278481871381   0.5575119762666707   0.4807751352808916   0.6478499859268729   0.9515080139328699   0.718976603594262   0.10920157180821849   0.838075530940331   0.8906999731612762   0.8786734987237037   0.805239485750448   0.889822815863025   0.46980966656267975   0.7515264951643491   0.5168923522216403   0.9448072902664494   0.13575505707605748   0.05986089386192219   0.7136769216195629   0.38521611081316703   0.6913908440676936   0.6760224118840628   0.9153280889817059   0.9795240784953702   0.11156299588055542   0.118510435617392   0.4345529537008143   0.33167409256849717   0.16005498194768555   0.39953383202313   0.3253513818925958   0.4935985616281661   0.2693550087864093   0.5208603332994263   0.5201118961421478   0.6037757457651411   0.7995453422237295   0.7693338381350772   0.0032195439205074793   0.6589684554986918   0.6637902851476721   0.709472944273155   0.28954262230094463   0.27375234468552473   0.9723994410799786   0.033450532389092236   0.37421453331923876
0.29422826619015463   0.8608364451994232   0.9149400967717002   0.9396615796184244   0.9625541736216574   0.7007814632517376   0.5154062647485702   0.6143101977258286   0.46895561199349134   0.4314264544653283   0.9945459314491439   0.0941983015836809   0.8651798662283502   0.6318811122415987   0.22521209331406683   0.09097875766317341   0.20621141072965846   0.9680908270939267   0.5157391490409119   0.8014361353622288   0.9324590660441338   0.995691386013948   0.48228861665181966   0.42722160204299003   0.6382307998539791   0.13485494081452493   0.5673485198801195   0.48756002242456553   0.6756766262323216   0.43407347756278736   0.05194225513154919   0.8732498246987369   0.20672101423883033   0.00264702309745903   0.057396323682405215   0.779051523115056   0.34154114801048013   0.3707659108558603   0.8321842303683383   0.6880727654518826   0.13532973728082165   0.40267508376193367   0.3164450813274265   0.8866366300896538   0.20287067123668795   0.4069836977479856   0.8341564646756068   0.4594150280466638   0.5646398713827089   0.2721287569334606   0.2668079447954874   0.9718550056220983   0.8889632451503872   0.8380552793706733   0.2148656896639382   0.09860518092336136   0.6822422309115569   0.8354082562732142   0.157469365981533   0.31955365780830536   0.3407010829010767   0.464642345417354   0.3252851356131946   0.6314808923564228
0.20537134562025505   0.06196726165542034   0.008840054285768131   0.744844262266769   0.002500674383567109   0.6549835639074347   0.1746835896101613   0.2854292342201052   0.4378608030008583   0.3828548069739741   0.9078756448146739   0.31357422859800693   0.5488975578504711   0.5447995276033009   0.6930099551507357   0.21496904767464559   0.8666553269389142   0.7093912713300865   0.5355405891692027   0.8954153898663403   0.5259542440378375   0.24474892591273256   0.2102554535560081   0.26393449750991743   0.32058289841758253   0.1827816642573122   0.20141539927023996   0.5190902352431485   0.31808222403401537   0.5277981003498774   0.02673180966007866   0.23366100102304327   0.8802214210331571   0.1449432933759033   0.11885616484540475   0.9200867724250363   0.33132386318268603   0.6001437657726025   0.425846209694669   0.7051177247503907   0.46466853624377175   0.8907524944425159   0.8903056205254664   0.8097023348840505   0.9387142922059342   0.6460035685297834   0.6800501669694582   0.545767837374133   0.6181313937883517   0.4632219042724712   0.47863476769921826   0.02667760213098458   0.30004916975433626   0.9354238039225937   0.4519029580391396   0.7930166011079413   0.4198277487211792   0.7904805105466904   0.3330467931937348   0.872929828682905   0.08850388553849316   0.1903367447740879   0.9072005834990658   0.16781210393251428
0.6238353492947214   0.299584250331572   0.016894962973599482   0.35810976904846376   0.6851210570887872   0.6535806818017886   0.33684479600414124   0.8123419316743308   0.06698966330043554   0.19035877752931743   0.858210028304923   0.7856643295433462   0.7669404935460993   0.2549349736067237   0.40630707026578344   0.9926477284354048   0.3471127448249201   0.4644544630600333   0.0732602770720486   0.11971789975249987   0.2586088592864269   0.2741177182859454   0.1660596935729828   0.9519057958199856   0.6347735099917055   0.9745334679543733   0.14916473059938332   0.5937960267715218   0.9496524529029183   0.3209527861525848   0.8123199345952421   0.7814540950971911   0.8826627896024828   0.1305940086232674   0.954109906290319   0.9957897655538449   0.1157222960563835   0.8756590350165436   0.5478028360245356   0.003142037118440069   0.7686095512314635   0.4112045719565104   0.474542558952487   0.8834241373659402   0.5100006919450365   0.13708685367056503   0.3084828653795042   0.9315183415459546   0.8752271819533309   0.16255338571619163   0.15931813478012088   0.33772231477443276   0.9255747290504127   0.8416005995636069   0.3469982001848788   0.5562682196772417   0.04291193944792997   0.7110065909403395   0.3928882938945598   0.5604784541233968   0.9271896433915465   0.8353475559237957   0.8450854578700242   0.5573364170049567
0.15858009216008306   0.4241429839672854   0.3705428989175372   0.6739122796390165   0.6485794002150466   0.28705613029672034   0.06206003353803302   0.7423939380930619   0.7733522182617155   0.12450274458052871   0.9027418987579121   0.4046716233186291   0.8477774892113029   0.28290214501692185   0.5557436985730333   0.8484034036413874   0.8048655497633729   0.5718955540765824   0.1628554046784735   0.28792494951799064   0.8776759063718265   0.7365479981527866   0.31776994680844933   0.7305885325130339   0.7190958142117434   0.31240501418550126   0.947227047890912   0.05667625287401742   0.07051641399669681   0.025348883888780916   0.885167014352879   0.31428231478095553   0.29716419573498126   0.9008461393082522   0.9824251155949669   0.9096106914623264   0.4493867065236784   0.6179439942913303   0.42668141702193363   0.06120728782093898   0.6445211567603055   0.04604844021474793   0.2638260123434601   0.7732823383029483   0.7668452503884791   0.3095004420619613   0.9460560655350108   0.04269380578991442   0.047749436176735674   0.99709542787646   0.9988290176440987   0.986017552915897   0.9772330221800388   0.9717465439876791   0.1136620032912196   0.6717352381349415   0.6800688264450576   0.0709004046794269   0.13123688769625266   0.7621245466726151   0.23068211992137924   0.4529564103880966   0.704555470674319   0.7009172588516761
0.5861609631610738   0.4069079701733486   0.4407294583308589   0.9276349205487278   0.8193157127725947   0.09740752811138734   0.49467339279584815   0.8849411147588133   0.7715662765958591   0.10031210023492731   0.49584437515174945   0.8989235618429163   0.7943332544158201   0.1285655562472482   0.38218237186052983   0.22718832370797484   0.11426442797076257   0.05766515156782129   0.2509454841642772   0.4650637770353597   0.8835823080493833   0.6047087411797247   0.5463900134899582   0.7641465181836836   0.29742134488830957   0.19780077100637608   0.10566055515909925   0.8365115976349559   0.47810563211571483   0.10039324289498874   0.6109871623632511   0.9515704828761425   0.7065393555198558   0.00008114266006143214   0.11514278721150166   0.052646921033226234   0.9122061011040355   0.8715155864128132   0.7329604153509718   0.8254585973252514   0.797941673133273   0.813850434844992   0.4820149311866946   0.3603948202898916   0.9143593650838897   0.20914169366526722   0.9356249176967364   0.5962483021062079   0.6169380201955802   0.011340922658891136   0.8299643625376372   0.7597367044712521   0.1388323880798653   0.9109476797639023   0.21897720017438607   0.8081662215951095   0.4322930325600095   0.9108665371038409   0.1038344129628844   0.7555193005618833   0.520086931455974   0.039350950691027724   0.3708739976119126   0.9300607032366319
0.7221452583227009   0.22550051584603578   0.888859066425218   0.5696658829467403   0.8077858932388112   0.01635882218076855   0.9532341487284816   0.9734175808405323   0.19084787304323103   0.0050178995218774156   0.12326978619084439   0.21368087636928018   0.052015484963365714   0.09407021975797503   0.9042925860164583   0.40551465477417065   0.6197224524033562   0.18320368265413406   0.8004581730535739   0.6499953542122874   0.09963552094738225   0.14385273196310633   0.42958417544166133   0.7199346509756555   0.3774902626246813   0.9183522161170705   0.5407251090164433   0.15026876802891517   0.5697043693858702   0.901993393936302   0.5874909602879618   0.17685118718838289   0.3788564963426391   0.8969754944144246   0.4642211740971174   0.9631703108191028   0.3268410113792734   0.8029052746564496   0.559928588080659   0.5576556560449321   0.7071185589759172   0.6197015920023156   0.7594704150270851   0.9076603018326448   0.607483038028535   0.4758488600392092   0.3298862395854238   0.1877256508569893   0.22999277540385363   0.5574966439221386   0.7891611305689804   0.03745688282807414   0.6602884060179834   0.6555032499858366   0.2016701702810187   0.8606056956396912   0.2814319096753443   0.7585277555714119   0.7374489961839014   0.8974353848205885   0.9545908982960709   0.9556224809149624   0.1775204081032423   0.3397797287756565
0.24747233932015367   0.33592088891264693   0.4180499930761572   0.43211942694301175   0.6399893012916187   0.8600720288734377   0.08816375349073341   0.24439377608602242   0.40999652588776503   0.30257538495129915   0.29900262292175295   0.20693689325794828   0.7497081198697816   0.6470721349654626   0.09733245264073428   0.34633119761825704   0.4682762101944372   0.8885443793940505   0.35988345645683295   0.4488958127976685   0.5136853118983663   0.9329218984790881   0.18236304835359066   0.10911608402201203   0.26621297257821264   0.5970010095664412   0.7643130552774334   0.6769966570790003   0.626223671286594   0.7369289806930035   0.6761493017867001   0.4326028809929779   0.21622714539882895   0.4343535957417043   0.37714667886494707   0.22566598773502958   0.4665190255290474   0.7872814607762417   0.2798142262242128   0.8793347901167725   0.9982428153346101   0.8987370813821912   0.9199307697673799   0.430438977319104   0.4845575034362438   0.9658151829031031   0.7375677214137892   0.321322893297092   0.21834453085803118   0.36881417333666183   0.9732546661363557   0.6443262362180917   0.5921208595714372   0.6318851926436584   0.2971053643496556   0.21172335522511385   0.37589371417260825   0.1975315969019541   0.9199586854847085   0.9860573674900842   0.9093746886435609   0.4102501361257123   0.6401444592604957   0.1067225773733117
0.9111318733089507   0.5115130547435212   0.7202136894931158   0.6762836000542076   0.42657436987270686   0.5456978718404181   0.9826459680793267   0.35496070675711566   0.20822983901467568   0.17688369850375618   0.009391301942970984   0.710634470539024   0.6161089794432385   0.5449985058600978   0.7122859375933154   0.4989111153139101   0.24021526527063025   0.3474669089581437   0.7923272521086068   0.5128537478238259   0.3308405766270694   0.9372167728324314   0.1521827928481111   0.40613117045051417   0.4197087033181187   0.4257037180889103   0.4319691033549952   0.7298475703963064   0.9931343334454118   0.8800058462484922   0.44932313527566853   0.3748868636391908   0.7849044944307362   0.703122147744736   0.43993183333269753   0.6642523931001669   0.16879551498749767   0.15812364188463823   0.7276458957393822   0.1653412777862568   0.9285802497168674   0.8106567329264945   0.9353186436307754   0.652487529962431   0.597739673089798   0.8734399600940631   0.7831358507826643   0.2463563595119168   0.17803096977167931   0.4477362420051529   0.35116674742766907   0.5165087891156104   0.1848966363262675   0.5677303957566606   0.9018436121520005   0.1416219254764195   0.39999214189553134   0.8646082480119246   0.461911778819303   0.47736953237625257   0.23119662690803366   0.7064846061272865   0.7342658830799208   0.3120282545899958
0.30261637719116624   0.8958278732007919   0.7989472394491454   0.6595407246275649   0.7048767041013683   0.022387913106728767   0.015811388666481102   0.413184365115648   0.5268457343296888   0.5746516711015759   0.6646446412388121   0.8966755760000377   0.3419490980034214   0.0069212753449152216   0.7628010290868115   0.7550536505236182   0.9419569561078901   0.14231302733299056   0.3008892502675085   0.2776841181473656   0.7107603291998564   0.43582842120570414   0.5666233671875878   0.9656558635573699   0.40814395200869014   0.5400005480049123   0.7676761277384423   0.306115138929805   0.703267247907322   0.5176126348981834   0.7518647390719613   0.892930773814157   0.17642151357763305   0.9429609637966075   0.0872200978331492   0.9962551978141193   0.8344724155742116   0.9360396884516924   0.3244190687463377   0.2412015472905011   0.8925154594663216   0.7937266611187018   0.023529818478829193   0.9635174291431354   0.18175513026646517   0.35789823991299763   0.45690645129124147   0.9978615655857657   0.773611178257775   0.8178976919080854   0.6892303235527991   0.6917464266559606   0.07034393035045308   0.30028505700990193   0.937365584480838   0.7988156528418037   0.89392241677282   0.35732409321329434   0.8501454866476887   0.8025604550276844   0.05945000119860838   0.42128440476160195   0.525726417901351   0.5613589077371832
0.1669345417322868   0.6275577436429002   0.5021965994225218   0.5978414785940478   0.9851794114658217   0.26965950372990255   0.04529014813128036   0.5999799130082821   0.21156823320804663   0.4517618118218171   0.35605982457848123   0.9082334863523215   0.14122430285759355   0.1514767548119152   0.4186942400976433   0.10941783351051784   0.24730188608477352   0.7941526615986209   0.5685487534499546   0.3068573784828335   0.18785188488616514   0.3728682568370189   0.04282233554860357   0.7454984707456502   0.020917343153878318   0.7453105131941187   0.5406257361260818   0.14765699215160252   0.03573793168805668   0.4756510094642162   0.4953355879948014   0.5476770791433204   0.8241696984800101   0.02388919764239908   0.13927576341632017   0.6394435927909989   0.6829453956224165   0.8724124428304839   0.7205815233186769   0.5300257592804811   0.435643509537643   0.07825978123186302   0.1520327698687223   0.2231683807976476   0.2477916246514779   0.7053915243948441   0.10921043432011872   0.4776699100519973   0.22687428149759956   0.9600810112007254   0.568584698194037   0.3300129179003948   0.19113634980954286   0.4844300017365092   0.07324911019923558   0.7823358387570744   0.3669666513295328   0.4605408040941101   0.9339733467829154   0.14289224596607542   0.6840212557071162   0.5881283612636262   0.21339182346423854   0.6128664866855943
0.24837774616947328   0.5098685800317632   0.06135905359551624   0.38969810588794673   0.0005861215179954072   0.8044770556369191   0.9521486192753975   0.9120281958359494   0.7737118400203958   0.8443960444361938   0.38356392108136056   0.5820152779355546   0.582575490210853   0.3599660426996845   0.310314810882125   0.7996794391784803   0.21560883888132015   0.8994252386055744   0.37634146409920954   0.6567871932124049   0.5315875831742038   0.31129687734194816   0.16294964063497103   0.043920706526810536   0.28320983700473057   0.801428297310185   0.10159058703945477   0.6542226006388638   0.2826237154867352   0.9969512416732659   0.14944196776405724   0.7421944048029143   0.5089118754663393   0.15255519723707217   0.7658780466826968   0.1601791268673597   0.9263363852554863   0.7925891545373877   0.4555632358005718   0.3604996876888794   0.7107275463741662   0.8931639159318132   0.07922177170136221   0.7037124944764745   0.1791399631999623   0.581867038589865   0.9162721310663912   0.659791787949664   0.8959301261952317   0.78043874127968   0.8146815440269364   0.0055691873108002065   0.6133064107084966   0.7834874996064142   0.6652395762628792   0.2633747825078859   0.10439453524215722   0.6309323023693421   0.8993615295801825   0.10319565564052617   0.17805814998667086   0.8383431478319544   0.4437982937796107   0.7426959679516467
0.46733060361250467   0.9451792319001411   0.3645765220782485   0.03898347347517224   0.28819064041254233   0.3633121933102761   0.44830439101185726   0.37919168552550825   0.3922605142173106   0.582873452030596   0.6336228469849209   0.37362249821470805   0.7789541035088141   0.7993859524241819   0.9683832707220417   0.11024771570682218   0.6745595682666569   0.16845365005483987   0.06902174114185922   0.007052060066296013   0.496501418279986   0.3301105022228855   0.6252234473622486   0.2643560921146492   0.029170814667481327   0.3849312703227444   0.2606469252840001   0.225372618639477   0.740980174254939   0.02161907701246826   0.8123425342721428   0.8461809331139688   0.34871966003762833   0.4387456249818722   0.17871968728722193   0.47255843489926075   0.5697655565288143   0.6393596725576903   0.21033641656518023   0.36231071919243857   0.8952059882621575   0.4709060225028505   0.14131467542332102   0.3552586591261425   0.39870456998217146   0.140795520279965   0.5160912280610725   0.0909025670114933   0.3695337553146901   0.7558642499572207   0.2554443027770724   0.8655299483720162   0.6285535810597511   0.7342451729447523   0.44310176850492966   0.01934901525804752   0.2798339210221228   0.2954995479628802   0.26438208121770773   0.5467905803587868   0.7100683644933085   0.6561398754051898   0.0540456646525275   0.18447986116634824
0.8148623762311511   0.18523385290233932   0.9127309892292065   0.8292212020402057   0.41615780624897963   0.04443833262237432   0.396639761168134   0.7383186350287124   0.04662405093428951   0.28857408266515366   0.14119545839106154   0.8727886866566962   0.4180704698745384   0.5543289097204013   0.6980936898861319   0.8534396713986486   0.1382365488524156   0.25882936175752114   0.4337116086684241   0.3066490910398618   0.4281681843591071   0.6026894863523313   0.37966594401589665   0.12216922987351357   0.613305808127956   0.417455633449992   0.46693495478669017   0.29294802783330787   0.1971480018789764   0.3730173008276177   0.07029519361855617   0.5546293928045954   0.1505239509446869   0.08444321816246399   0.9290997352274947   0.6818407061478993   0.7324534810701485   0.5301143084420626   0.23100604534136276   0.8284010347492508   0.594216932217733   0.27128494668454156   0.7972944366729386   0.5217519437093889   0.16604874785862586   0.6685954603322102   0.417628492657042   0.39958271383587535   0.5527429397306698   0.25113982688221825   0.9506935378703518   0.10663468600256748   0.35559493785169344   0.8781225260546006   0.8803983442517956   0.552005293197972   0.2050709869070065   0.7936793078921366   0.9512986090243011   0.8701645870500727   0.47261750583685797   0.2635649994500739   0.7202925636829383   0.041763552300822016
0.878400573619125   0.9922800527655323   0.9229981270099997   0.5200116085914331   0.7123518257604992   0.3236845924333221   0.5053696343529577   0.12042889475555779   0.1596088860298293   0.07254476555110388   0.5546760964826059   0.01379420875299031   0.8040139481781359   0.1944222394965033   0.6742777522308101   0.4617889155550183   0.5989429612711294   0.40074293160436675   0.7229791432065091   0.5916243285049455   0.12632545543427143   0.13717793215429283   0.0026865795235707793   0.5498607762041235   0.24792488181514644   0.14489787938876048   0.0796884525135711   0.02984916761269042   0.5355730560546473   0.8212132869554384   0.5743188181606134   0.9094202728571327   0.37596417002481797   0.7486685214043345   0.019642721678007586   0.8956260641041424   0.5719502218466821   0.5542462819078312   0.34536496944719747   0.43383714854912403   0.9730072605755526   0.15350335030346446   0.6223858262406884   0.8422128200441785   0.8466818051412812   0.01632541814917163   0.6196992467171176   0.292352043840055   0.5987569233261348   0.8714275387604111   0.5400107942035465   0.2625028762273645   0.06318386727148753   0.05021425180497277   0.9656919760429331   0.3530826033702319   0.6872196972466695   0.30154573040063826   0.9460492543649255   0.4574565392660896   0.1152694753999875   0.747299448492807   0.6006842849177281   0.02361939071696553
0.14226221482443482   0.5937960981893426   0.9782984586770397   0.18140657067278704   0.2955804096831536   0.577470680040171   0.3585992119599221   0.8890545268327321   0.6968234863570187   0.7060431412797599   0.8185884177563756   0.6265516506053675   0.6336396190855312   0.6558288894747871   0.8528964417134426   0.27346904723513565   0.9464199218388617   0.3542831590741488   0.9068471873485171   0.816012507969046   0.8311504464388741   0.6069837105813417   0.3061629024307891   0.7923931172520805   0.6888882316144394   0.013187612391999096   0.3278644437537494   0.6109865465792935   0.3933078219312858   0.4357169323518281   0.9692652317938273   0.7219320197465614   0.696484335574267   0.7296737910720683   0.15067681403745165   0.09538036914119387   0.0628447164887358   0.07384490159728119   0.2977803723240091   0.8219113219060582   0.11642479464987414   0.7195617425231324   0.390933184975492   0.005898813937012174   0.28527434821099995   0.11257803194179068   0.08477028254470292   0.21350569668493163   0.5963861165965606   0.09939041954979158   0.7569058387909535   0.6025191501056382   0.20307829466527483   0.6636734871979635   0.7876406069971262   0.8805871303590768   0.5065939590910078   0.9339996961258952   0.6369637929596746   0.7852067612178829   0.443749242602272   0.860154794528614   0.33918342063566553   0.9632954393118246
0.32732444795239785   0.14059305200548164   0.9482502356601735   0.9573966253748124   0.0420500997413979   0.02801502006369095   0.8634799531154707   0.7438909286898808   0.4456639831448373   0.9286246005138994   0.10657411432451705   0.14137177858424266   0.2425856884795625   0.2649511133159359   0.3189335073273908   0.26078464822516595   0.7359917293885547   0.3309514171900407   0.6819697143677161   0.47557788700728304   0.29224248678628273   0.4707966226614267   0.34278629373205066   0.5122824476954585   0.9649180388338848   0.330203570655945   0.39453605807187714   0.554885822320646   0.922867939092487   0.3021885505922541   0.5310561049564065   0.8109948936307652   0.47720395594764964   0.37356395007835475   0.42448199063188946   0.6696231150465225   0.23461826746808714   0.10861283676241883   0.10554848330449867   0.4088384668213566   0.49862653807953244   0.7776614195723781   0.4235787689367825   0.9332605798140735   0.20638405129324974   0.3068647969109515   0.08079247520473185   0.4209781321186151   0.24146601245936491   0.9766612262550064   0.6862564171328547   0.8660923097979691   0.31859807336687795   0.6744726756627524   0.1552003121764482   0.055097416167203914   0.8413941174192283   0.30090872558439763   0.7307183215445587   0.3854743011206814   0.6067758499511412   0.1922958888219788   0.6251698382400601   0.9766358342993248
0.10814931187160874   0.4146344692496006   0.20159106930327758   0.04337525448525122   0.901765260578359   0.10776967233864918   0.12079859409854574   0.6223971223666361   0.6602992481189941   0.13110844608364275   0.43454217696569103   0.756304812568667   0.3417011747521161   0.4566357704208904   0.27934186478924283   0.7012073964014631   0.5003070573328877   0.15572704483649277   0.5486235432446841   0.3157330952807817   0.8935312073817466   0.963431156014514   0.923453705004624   0.3390972609814569   0.7853818955101378   0.5487966867649133   0.7218626357013465   0.2957220064962057   0.8836166349317789   0.4410270144262642   0.6010640416028007   0.6733248841295696   0.22331738681278476   0.30991856834262144   0.1665218646371097   0.9170200715609026   0.8816162120606686   0.853282797921731   0.8871799998478669   0.2158126751594395   0.38130915472778093   0.6975557530852382   0.3385564566031828   0.9000795798786577   0.4877779473460343   0.7341245970707243   0.41510275159855875   0.5609823188972008   0.7023960518358965   0.18532791030581094   0.6932401158972124   0.26526031240099507   0.8187794169041176   0.7443008958795467   0.09217607429441162   0.5919354282714255   0.5954620300913329   0.43438232753692535   0.9256542096573019   0.6749153567105229   0.7138458180306642   0.5810995296151943   0.03847420980943505   0.4591026815510834
0.3325366633028833   0.8835437765299561   0.6999177532062523   0.5590231016724256   0.8447587159568489   0.1494191794592318   0.28481500160769346   0.9980407827752248   0.14236266412095247   0.9640912691534209   0.5915748857104811   0.7327804703742298   0.32358324721683485   0.2197903732738741   0.4993988114160695   0.14084504210280424   0.7281212171255019   0.7854080457369488   0.5737446017587676   0.46592968539228136   0.014275399094837781   0.20430851612175444   0.5352703919493326   0.0068270038411979445   0.6817387357919545   0.32076473959179835   0.8353526387430803   0.4478039021687723   0.8369800198351055   0.17134556013256655   0.5505376371353868   0.4497631193935475   0.6946173557141531   0.20725429097914566   0.9589627514249057   0.7169826490193177   0.3710341084973182   0.9874639177052715   0.45956394000883616   0.5761376069165135   0.6429128913718163   0.2020558719683228   0.8858193382500685   0.11020792152423219   0.6286374922769785   0.9977473558465684   0.350548946300736   0.10338091768303424   0.946898756485024   0.6769826162547701   0.5151963075576557   0.655577015514262   0.10991873664991846   0.5056370561222034   0.9646586704222689   0.20581389612071443   0.4153013809357654   0.2983827651430578   0.005695918997363212   0.48883124710139664   0.044267272438447164   0.31091884743778625   0.5461319789885271   0.9126936401848831
0.4013543810666309   0.10886297546946343   0.6603126407384585   0.8024857186606509   0.7727168887896524   0.11111561962289505   0.3097636944377225   0.6991048009776167   0.8258181323046284   0.43413300336812505   0.7945673868800668   0.04352778546335476   0.7158993956547101   0.9284959472459215   0.829908716457798   0.8377138893426403   0.3005980147189446   0.6301131821028637   0.8242127974604347   0.34888264224124366   0.25633074228049746   0.3191943346650775   0.27808081847190763   0.4361890020563605   0.8549763612138666   0.21033135919561408   0.6177681777334492   0.6337032833957096   0.08225947242421411   0.09921573957271901   0.3080044832957266   0.934598482418093   0.25644134011958564   0.665082736204594   0.5134370964156598   0.8910706969547382   0.5405419444648757   0.7365867889586725   0.683528379957862   0.053356807612097844   0.23994392974593104   0.10647360685580871   0.8593155824974272   0.7044741653708542   0.9836131874654336   0.7872792721907312   0.5812347640255195   0.26828516331449365   0.12863682625156705   0.5769479129951172   0.9634665862920705   0.634581879918784   0.04637735382735293   0.47773217342239815   0.6554621029963439   0.699983397500691   0.7899360137077672   0.8126494372178041   0.142025006580684   0.8089127005459529   0.24939406924289162   0.0760626482591317   0.4584966266228221   0.7555558929338551
0.00945013949696058   0.969589041403323   0.5991810441253949   0.05108172756300091   0.025836952031526993   0.1823097692125918   0.01794628009987526   0.7827965642485073   0.89720012577996   0.6053618562174746   0.05447969380780479   0.14821468432972326   0.850822771952607   0.1276296827950765   0.39901759081146093   0.4482312868290322   0.06088675824483975   0.31498024557727233   0.2569925842307769   0.6393185862830792   0.8114926890019482   0.23891759731814063   0.7984959576079549   0.8837626933492242   0.8020425495049875   0.26932855591481764   0.19931491348256   0.8326809657862233   0.7762055974734605   0.08701878670222586   0.18136863338268475   0.04988440153771598   0.8790054716935006   0.4816569304847512   0.12688893957487996   0.9016697172079927   0.02818269974089358   0.35402724768967475   0.727871348763419   0.45343843037896053   0.9672959414960538   0.03904700211240239   0.47087876453264205   0.8141198440958812   0.1558032524941057   0.8001294047942618   0.6723828069246872   0.9303571507466571   0.35376070298911816   0.5308008488794441   0.4730678934421272   0.09767618496043384   0.5775551055156576   0.4437820621772183   0.29169926005944247   0.047791783422717865   0.698549633822157   0.962125131692467   0.1648103204845625   0.14612206621472515   0.6703669340812634   0.6080978840027923   0.43693897172114354   0.6926836358357646
0.7030709925852096   0.5690508818903899   0.9660602071885015   0.8785637917398834   0.5472677400911039   0.7689214770961281   0.2936774002638143   0.9482066409932263   0.19350703710198572   0.23812062821668403   0.8206095068216871   0.8505304560327924   0.6159519315863281   0.7943385660394658   0.5289102467622446   0.8027386726100746   0.9174022977641711   0.8322134343469988   0.3640999262776821   0.6566166063953494   0.24703536368290774   0.2241155503442065   0.9271609545565386   0.9639329705595847   0.5439643710976981   0.6550646684538166   0.9611007473680371   0.08536917881970141   0.9966966310065943   0.8861431913576885   0.6674233471042228   0.13716253782647514   0.8031895939046085   0.6480225631410044   0.8468138402825357   0.2866320817936827   0.1872376623182804   0.8536839971015386   0.31790359352029113   0.4838934091836082   0.2698353645541093   0.021470562754539825   0.953803667242609   0.8272768027882588   0.02280000087120152   0.7973550124103334   0.026642712686070456   0.863343832228674   0.47883562977350336   0.14229034395651674   0.06554196531803337   0.7779746534089725   0.4821389987669091   0.2561471525988283   0.39811861821381056   0.6408121155824975   0.6789494048623005   0.6081245894578239   0.5513047779312749   0.35418003378881474   0.4917117425440201   0.7544405923562852   0.2334011844109837   0.8702866246052066
0.22187637798991086   0.7329700296017454   0.27959751716837467   0.043009821816947826   0.19907637711870935   0.9356150171914122   0.25295480448230423   0.17966598958827384   0.7202407473452059   0.7933246732348954   0.18741283916427087   0.40169133617930125   0.2381017485782969   0.537177520636067   0.7892942209504603   0.7608792205968038   0.5591523437159964   0.9290529311782432   0.23798944301918548   0.40669918680798905   0.06744060117197626   0.17461233882195795   0.004588258608201784   0.5364125622027824   0.8455642231820654   0.44164230922021247   0.7249907414398271   0.49340274038583465   0.6464878460633561   0.5060272920288004   0.4720359369575229   0.3137367507975608   0.9262470987181501   0.712702618793905   0.284623097793252   0.9120454146182596   0.6881453501398532   0.1755250981578379   0.4953288768427917   0.15116619402145579   0.1289930064238568   0.24647216697959468   0.2573394338236062   0.7444670072134667   0.06155240525188056   0.07185982815763674   0.2527511752154044   0.20805444501068426   0.21598818206981515   0.6302175189374243   0.5277604337755774   0.7146517046248496   0.5695003360064591   0.12419022690862386   0.055724496818054456   0.4009149538272888   0.643253237288309   0.41148760811471885   0.7711013990248025   0.48886953920902926   0.9551078871484558   0.23596250995688095   0.27577252218201076   0.3377033451875735
0.826114880724599   0.9894903429772863   0.018433088358404535   0.5932363379741068   0.7645624754727184   0.9176305148196495   0.7656819131430002   0.3851818929634225   0.5485742934029033   0.2874129958822253   0.23792147936742278   0.6705301883385728   0.9790739573964442   0.16322276897360144   0.18219698254936834   0.269615234511284   0.3358207201081352   0.7517351608588826   0.4110955835245659   0.7807456953022547   0.3807128329596794   0.5157726509020016   0.13532306134255515   0.44304235011468124   0.5545979522350803   0.5262823079247153   0.1168899729841506   0.8498060121405745   0.790035476762362   0.6086517931050658   0.3512080598411505   0.464624119177152   0.24146118335945865   0.3212387972228405   0.11328658047372771   0.7940939308385792   0.26238722596301445   0.15801602824923905   0.9310895979243594   0.5244786963272952   0.9265665058548793   0.40628086739035646   0.5199940143997935   0.7437330010250405   0.5458536728951999   0.8905082164883549   0.38467095305723836   0.3006906509103592   0.9912557206601196   0.3642259085636395   0.26778098007308776   0.4508846387697847   0.20122024389775764   0.7555741154585737   0.9165729202319373   0.9862605195926327   0.959759060538299   0.43433531823573324   0.8032863397582095   0.1921665887540535   0.6973718345752845   0.2763192899864942   0.8721967418338502   0.6676878924267583
0.7708053287204052   0.8700384225961377   0.3522027274340567   0.9239548914017179   0.2249516558252053   0.9795302061077829   0.9675317743768183   0.6232642404913588   0.23369593516508574   0.6153042975441433   0.6997507943037306   0.17237960172157404   0.03247569126732811   0.8597301820855696   0.7831778740717933   0.18611908212894135   0.07271663072902913   0.4253948638498364   0.9798915343135838   0.9939524933748879   0.3753447961537446   0.14907557386334222   0.10769479247973363   0.3262646009481295   0.6045394674333394   0.2790371512672045   0.755492065045677   0.4023097095464116   0.3795878116081341   0.29950694515942167   0.7879602906688586   0.7790454690550529   0.14589187644304838   0.6842026476152784   0.08820949636512809   0.6066658673334788   0.11341618517572026   0.8244724655297087   0.3050316222933348   0.4205467852045375   0.04069955444669113   0.39907760167987233   0.325140087979751   0.4265942918296496   0.6653547582929465   0.2500020278165301   0.21744529550001737   0.1003296908815201   0.06081529085960708   0.9709648765493256   0.46195323045434045   0.6980199813351086   0.681227479251473   0.6714579313899038   0.6739929397854818   0.9189745122800557   0.5353356028084246   0.9872552837746256   0.5857834434203537   0.31230864494657684   0.4219194176327043   0.16278281824491686   0.2807518211270189   0.8917618597420394
0.3812198631860132   0.7637052165650445   0.9556117331472679   0.4651675679123898   0.7158651048930667   0.5137031887485145   0.7381664376472505   0.3648378770308697   0.6550498140334596   0.5427383121991889   0.2762132071929101   0.6668178956957611   0.9738223347819867   0.871280380809285   0.6022202674074283   0.7478433834157054   0.4384867319735621   0.8840250970346595   0.01643682398707464   0.4355347384691286   0.01656731434085775   0.7212422787897426   0.7356850028600558   0.5437728787270892   0.6353474511548446   0.957537062224698   0.7800732697127878   0.07860531081469942   0.9194823462617778   0.4438338734761836   0.04190683206553729   0.7137674337838298   0.26443253222831825   0.9010955612769946   0.7656936248726272   0.046949538088068565   0.2906101974463316   0.02981518046770968   0.16347335746519887   0.29910615467236307   0.8521234654727695   0.14579008343305025   0.14703653347812423   0.8635714162032344   0.8355561511319118   0.42454780464330766   0.4113515306180685   0.31979853747614523   0.20020869997706722   0.4670107424186096   0.6312782609052807   0.2411932266614458   0.28072635371528937   0.023176868942426043   0.5893714288397434   0.527425792877616   0.016293821486971092   0.12208130766543136   0.8236778039671162   0.48047625478954753   0.7256836240406395   0.09226612719772168   0.6602044465019173   0.18137010011718444
0.87356015856787   0.9464760437646714   0.5131679130237932   0.31779868391395   0.03800400743595816   0.5219282391213638   0.10181638240572463   0.9980001464378048   0.837795307458891   0.05491749670275416   0.47053812150044394   0.7568069197763589   0.5570689537436015   0.03174062776032811   0.8811666926607006   0.22938112689874288   0.5407751322566305   0.9096593200948968   0.057488888693584365   0.7489048721091953   0.815091508215991   0.817393192897175   0.39728444219166703   0.567534771992011   0.941531349648121   0.8709171491325036   0.8841165291678739   0.24973608807806097   0.9035273422121629   0.34898891001113985   0.7823001467621493   0.2517359416402562   0.06573203475327197   0.2940714133083857   0.3117620252617053   0.49492902186389726   0.5086630810096704   0.2623307855480576   0.43059533260100474   0.2655478949651544   0.9678879487530399   0.35267146545316086   0.37310644390742037   0.516643022855959   0.15279644053704888   0.5352782725559858   0.9758220017157534   0.9491082508639481   0.2112650908889278   0.6643611234234821   0.09170547254787946   0.6993721627858871   0.3077377486767649   0.3153722134123423   0.30940532578573016   0.4476362211456309   0.24200571392349296   0.021300800103956574   0.9976433005240248   0.9527071992817336   0.7333426329138226   0.758970014555899   0.5670479679230201   0.6871593043165792
0.7654546841607827   0.40629854910273816   0.1939415240155997   0.17051628146062026   0.6126582436237338   0.8710202765467524   0.21811952229984632   0.2214080305966722   0.40139315273480597   0.20665915312327027   0.12641404975196688   0.522035867810785   0.09365540405804107   0.891286939710928   0.8170087239662367   0.07439964666515417   0.8516496901345482   0.8699861396069715   0.8193654234422119   0.12169244738342051   0.11830705722072554   0.11101612505107242   0.25231745551919177   0.43453314306684127   0.3528523730599428   0.7047175759483343   0.05837593150359205   0.26401686160622095   0.740194129436209   0.8336972994015819   0.8402564092037457   0.04260883100954879   0.3388009767014031   0.6270381462783117   0.7138423594517789   0.5205729631987637   0.24514557264336198   0.7357512065673836   0.8968336354855422   0.44617331653360953   0.3934958825088139   0.8657650669604122   0.07746821204333032   0.32448086915018903   0.27518882528808836   0.7547489419093398   0.8251507565241386   0.8899477260833478   0.9223364522281455   0.05003136596100552   0.7667748250205465   0.6259308644771269   0.18214232279193646   0.21633406655942364   0.9265184158168008   0.583322033467578   0.8433413460905334   0.589295920281112   0.21267605636502196   0.06274907026881432   0.5981957734471713   0.8535447137137284   0.3158424208794798   0.6165757537352048
0.2046998909383575   0.9877796467533162   0.2383742088361495   0.2920948845850157   0.9295110656502692   0.2330307048439764   0.4132234523120109   0.40214715850166793   0.007174613422123678   0.18299933888297087   0.6464486272914644   0.7762162940245411   0.8250322906301872   0.9666652723235473   0.7199302114746635   0.19289426055696304   0.9816909445396539   0.3773693520424352   0.5072541551096416   0.13014519028814872   0.38349517109248243   0.5238246383287068   0.19141173423016178   0.513569436552944   0.17879528015412494   0.5360449915753907   0.9530375253940123   0.22147455196792826   0.2492842145038558   0.30301428673141423   0.5398140730820014   0.8193273934662604   0.2421096010817321   0.12001494784844334   0.893365445790537   0.04311109944171926   0.4170773104515449   0.15334967552489612   0.1734352343158735   0.8502168388847562   0.435386365911891   0.7759803234824609   0.6661810792062319   0.7200716485966074   0.051891194819408556   0.2521556851537541   0.47476934497607015   0.2065022120436635   0.8730959146652836   0.7161106935783634   0.5217318195820578   0.9850276600757353   0.6238117001614278   0.41309640684694926   0.9819177465000565   0.16570026660947493   0.3817020990796957   0.2930814589985059   0.0885523007095194   0.12258916716775568   0.9646247886281508   0.1397317834736098   0.9151170663936459   0.27237232828299945
0.5292384227162599   0.3637514599911489   0.248935987187414   0.552300679686392   0.4773472278968513   0.11159577483739479   0.7741666422113439   0.3457984676427285   0.6042513132315677   0.3954850812590313   0.252434822629286   0.3607708075669932   0.9804396130701398   0.982388674412082   0.2705170761292296   0.19507054095751825   0.5987375139904442   0.6893072154135761   0.18196477541971018   0.07248137378976258   0.6341127253622932   0.5495754319399663   0.26684770902606425   0.8001090455067631   0.10487430264603342   0.18582397194881745   0.017911721838650252   0.24780836582037113   0.6275270747491821   0.07422819711142264   0.24374507962730638   0.9020098981776427   0.02327576151761446   0.6787431158523913   0.9913102569980203   0.5412390906106495   0.04283614844747462   0.6963544414403093   0.7207931808687907   0.3461685496531312   0.4440986344570305   0.007047226026733167   0.5388284054490806   0.27368717586336866   0.8099859090947372   0.45747179408676686   0.2719806964230163   0.4735781303566055   0.7051116064487039   0.2716478221379494   0.25406897458436606   0.2257697645362344   0.07758453169952169   0.19741962502652677   0.010323894957059682   0.3237598663585917   0.05430877018190723   0.5186765091741354   0.019013637959039337   0.7825207757479423   0.01147262173443261   0.8223220677338261   0.2982204570902486   0.43635222609481106
0.5673739872774021   0.815274841707093   0.759392051641168   0.16266505023144243   0.7573880781826648   0.3578030476203261   0.4874113552181517   0.689086919874837   0.052276471733961036   0.08615522548237671   0.23334238063378565   0.4633171553386025   0.9746919400344394   0.88873560045585   0.22301848567672597   0.13955728898001077   0.9203831698525321   0.37005909128171455   0.20400484771768662   0.3570365132320685   0.9089105481180995   0.5477370235478884   0.905784390627438   0.9206842871372575   0.3415365608406974   0.7324621818407955   0.14639233898627002   0.758019236905815   0.5841484826580325   0.3746591342204693   0.6589809837681183   0.06893231703097809   0.5318720109240715   0.2885039087380926   0.42563860313433266   0.6056151616923756   0.5571800708896322   0.39976830828224263   0.20262011745760672   0.4660578727123648   0.6367969010371001   0.029709217000528126   0.9986152697399201   0.10902135948029634   0.7278863529190005   0.48197219345263975   0.09283087911248204   0.18833707234303892   0.3863497920783031   0.7495100116118443   0.946438540126212   0.4303178354372239   0.8022013094202706   0.37485087739137496   0.2874575563580937   0.36138551840624583   0.2703292984961991   0.08634696865328237   0.861818953223761   0.7557703567138703   0.713149227606567   0.6865786603710398   0.6591988357661543   0.2897124840015054
0.07635232656946692   0.6568694433705116   0.6605835660262342   0.18069112452120906   0.3484659736504664   0.17489724991787187   0.5677526869137521   0.9923540521781702   0.9621161815721633   0.4253872383060276   0.6213141467875402   0.5620362167409463   0.15991487215189268   0.0505363609146526   0.33385659042944643   0.20065069833470042   0.8895855736556936   0.9641893922613702   0.4720376372056854   0.4448803416208302   0.1764363460491266   0.27761073189033053   0.8128388014395311   0.15516785761932478   0.1000840194796597   0.6207412885198189   0.1522552354132969   0.9744767330981157   0.7516180458291933   0.44584403860194705   0.5845025484995447   0.9821226809199456   0.7895018642570301   0.0204568002959195   0.9631884017120046   0.4200864641789993   0.6295869921051374   0.9699204393812669   0.6293318112825581   0.21943576584429889   0.7400014184494438   0.005731047119896671   0.1572941740768727   0.7745554242234687   0.5635650724003172   0.7281203152295661   0.3444553726373416   0.619387566604144   0.4634810529206575   0.10737902670974722   0.1922001372240447   0.6449108335060282   0.7118630070914642   0.6615349881078002   0.6076975887245   0.6627881525860827   0.9223611428344342   0.6410781878118806   0.6445091870124954   0.2427016884070834   0.29277415072929674   0.6711577484306137   0.01517737572993721   0.023265922562784497
0.5527727322798529   0.6654267013107171   0.8578832016530645   0.2487104983393158   0.9892076598795357   0.9373063860811509   0.5134278290157229   0.6293229317351718   0.5257266069588783   0.8299273593714037   0.3212276917916782   0.9844120982291437   0.8138635998674141   0.16839237126360354   0.7135301030671782   0.32162394564306096   0.8915024570329799   0.5273141834517229   0.0690209160546829   0.07892225723597757   0.5987283063036832   0.8561564350211092   0.053843540324745684   0.055656334673193066   0.045955574023830256   0.19072973371039206   0.1959603386716812   0.8069458363338773   0.0567479141442945   0.2534233476292411   0.6825325096559584   0.17762290459870542   0.5310213071854162   0.4234959882578374   0.3613048178642801   0.19321080636956178   0.7171577073180021   0.2551036169942339   0.6477747147971018   0.8715868607265008   0.8256552502850222   0.727789433542511   0.578753798742419   0.7926646034905233   0.22692694398133897   0.8716329985214019   0.5249102584176732   0.7370082688173302   0.1809713699575087   0.6809032648110098   0.3289499197459921   0.9300624324834529   0.12422345581321421   0.42747991718176864   0.6464174100900337   0.7524395278847475   0.593202148627798   0.003983928923931212   0.2851125922257537   0.5592287215151858   0.8760444413097959   0.7488803119296973   0.6373378774286518   0.6876418607886849
0.05038919102477367   0.021090878387186335   0.05858407868623287   0.8949772572981617   0.8234622470434347   0.1494578798657845   0.5336738202685596   0.15796898848083143   0.642490877085926   0.4685546150547747   0.2047239005225675   0.22790655599737852   0.5182674212727117   0.041074697873006064   0.5583064904325338   0.47546702811263103   0.9250652726449138   0.03709076894907485   0.2731938982067801   0.9162383065974453   0.04902083133511794   0.28821045701937753   0.6358560207781282   0.22859644580876037   0.9986316403103442   0.2671195786321912   0.5772719420918954   0.33361918851059874   0.17516939326690958   0.1176616987664067   0.04359812182333577   0.17565020002976728   0.5326785161809836   0.649107083711632   0.8388742213007683   0.9477436440323888   0.014411094908271822   0.608032385838626   0.2805677308682345   0.4722766159197578   0.08934582226335804   0.570941616889551   0.0073738326614544636   0.5560383093223125   0.040324990928240094   0.28273115987017355   0.3715178118833262   0.32744186351355214   0.04169335061789582   0.015611581237982373   0.7942458697914309   0.9938226750029534   0.8665239573509862   0.8979498824715757   0.7506477479680951   0.8181724749731861   0.33384544117000264   0.2488427987599437   0.9117735266673268   0.8704288309407974   0.31943434626173084   0.6408104129213178   0.6312057957990923   0.3981522150210396
0.2300885239983728   0.06986879603176668   0.6238319631376379   0.8421139056987271   0.1897635330701327   0.7871376361615932   0.2523141512543116   0.5146720421851749   0.14807018245223688   0.7715260549236107   0.45806828146288076   0.5208493671822215   0.28154622510125066   0.8735761724520351   0.7074205334947856   0.7026768922090354   0.947700783931248   0.6247333736920914   0.7956470068274588   0.832248061268238   0.6282664376695172   0.9839229607707737   0.1644412110283665   0.4340958462471985   0.39817791367114436   0.9140541647390069   0.5406092478907286   0.5919819405484714   0.20841438060101167   0.12691652857741384   0.28829509663641706   0.07730989836329646   0.060344198148774786   0.3553904736538031   0.8302268151735362   0.5564605311810749   0.7787979730475242   0.481814301201768   0.12280628167875063   0.8537836389720395   0.8310971891162762   0.8570809275096767   0.3271592748512918   0.021535577703801406   0.202830751446759   0.873157966738903   0.1627180638229253   0.5874397314566029   0.8046528377756146   0.9591038019998961   0.6221088159321966   0.9954577909081315   0.596238457174603   0.8321872734224822   0.3338137192957796   0.9181478925448351   0.5358942590258282   0.47679679976867917   0.5035869041222433   0.3616873613637601   0.757096285978304   0.9949824985669111   0.38078062244349264   0.5079037223917207
0.9259990968620279   0.1379015710572345   0.05362134759220085   0.4863681446879192   0.7231683454152689   0.2647436043183315   0.8909032837692755   0.8989284132313163   0.9185155076396543   0.3056398023184354   0.26879446783707894   0.9034706223231849   0.3222770504650513   0.4734525288959532   0.9349807485412993   0.9853227297783498   0.7863827914392231   0.9966557291272741   0.43139384441905604   0.6236353684145897   0.029286505460919043   0.0016732305603629287   0.05061322197556339   0.11573164602286902   0.10328740859889116   0.8637716595031284   0.9969918743833626   0.6293635013349498   0.38011906318362226   0.599028055184797   0.10608859061408699   0.7304350881036334   0.46160355554396804   0.2933882528663615   0.8372941227770081   0.8269644657804486   0.13932650507891678   0.8199357239704084   0.9023133742357087   0.8416417360020988   0.3529437136396937   0.8232799948431343   0.4709195298166527   0.21800636758750916   0.32365720817877464   0.8216067642827714   0.4203063078410893   0.10227472156464014   0.22036979957988348   0.9578351047796428   0.42331443345772674   0.47291122022969034   0.8402507363962612   0.35880704959484594   0.31722584284363975   0.7424761321260569   0.37864718085229315   0.06541879672848444   0.4799317200666317   0.9155116663456083   0.2393206757733764   0.24548307275807613   0.577618345830923   0.0738699303435095
0.8863769621336827   0.4222030779149419   0.10669881601427031   0.8558635627560003   0.562719753954908   0.6005963136321706   0.686392508173181   0.7535888411913602   0.3423499543750246   0.6427612088525276   0.2630780747154543   0.2806776209616698   0.5020992179787634   0.2839541592576817   0.9458522318718146   0.5382014888356129   0.12345203712647025   0.21853536252919725   0.46592051180518285   0.6226898224900046   0.8841313613530939   0.9730522897711211   0.8883021659742598   0.5488198921464951   0.9977543992194111   0.5508492118561793   0.7816033499599895   0.6929563293904948   0.4350346452645031   0.9502528982240087   0.0952108417868085   0.9393674881991345   0.09268469088947849   0.3074916893714811   0.8321327670713542   0.6586898672374647   0.5905854729107151   0.023537530113799405   0.8862805351995396   0.12048837840185184   0.4671334357842448   0.8050021675846022   0.42036002339435685   0.49779855591184724   0.5830020744311509   0.8319498778134811   0.532057857420097   0.9489786637653521   0.5852476752117398   0.28110066595730177   0.7504545074601074   0.2560223343748574   0.15021302994723673   0.330847767733293   0.655243665673299   0.3166548461757228   0.057528339057758254   0.023356078361811923   0.8231108986019448   0.6579649789382581   0.46694286614704317   0.9998185482480125   0.9368303634024051   0.5374766005364062
0.9998094303627983   0.19481638066341037   0.5164703400080483   0.03967804462455899   0.41680735593164736   0.36286650284992933   0.9844124825879512   0.09069938085920685   0.8315596807199075   0.08176583689262759   0.23395797512784378   0.8346770464843495   0.6813466507726708   0.7509180691593346   0.5787143094545448   0.5180222003086267   0.6238183117149125   0.7275619907975227   0.7556034108526001   0.8600572213703686   0.15687544556786936   0.7277434425495102   0.818773047450195   0.3225806208339624   0.15706601520507102   0.5329270618860997   0.30230270744214666   0.28290257620940334   0.7402586592734237   0.17006055903617043   0.31789022485419544   0.19220319535019653   0.9086989785535161   0.08829472214354284   0.08393224972635166   0.35752614886584705   0.22735232778084535   0.33737665298420827   0.5052179402718069   0.8395039485572204   0.6035340160659328   0.6098146621866856   0.7496145294192068   0.9794467271868518   0.44665857049806346   0.8820712196371755   0.930841481969012   0.6568661063528894   0.28959255529299244   0.3491441577510757   0.6285387745268652   0.37396353014348604   0.5493338960195687   0.17908359871490528   0.3106485496726698   0.18176033479328954   0.6406349174660526   0.09078887657136243   0.22671629994631814   0.8242341859274425   0.41328258968520726   0.7534122235871542   0.7214983596745113   0.9847302373702221
0.8097485736192744   0.1435975614004686   0.9718838302553044   0.005283510183370319   0.363090003121211   0.2615263417632931   0.04104234828629255   0.34841740383048087   0.07349744782821854   0.9123821840122174   0.4125035737594273   0.9744538736869949   0.5241635518086498   0.7332985852973122   0.1018550240867575   0.7926935388937053   0.8835286343425972   0.6425097087259497   0.8751387241404394   0.9684593529662628   0.47024604465738995   0.8890974851387955   0.15364036446592808   0.9837291155960407   0.6604974710381155   0.745499923738327   0.18175653421062363   0.9784456054126703   0.29740746791690453   0.4839735819750338   0.14071418592433108   0.6300282015821895   0.22391002008868602   0.5715913979628164   0.7282106121649038   0.6555743278951947   0.6997464682800362   0.8382928126655043   0.6263555880781463   0.8628807890014893   0.8162178339374391   0.1957831039395546   0.7512168639377069   0.8944214360352265   0.34597178928004907   0.30668561880075906   0.5975764994717788   0.9106923204391858   0.6854743182419336   0.5611856950624322   0.41581996526115517   0.9322467150265155   0.388066850325029   0.07721211308739834   0.2751057793368241   0.302218513444326   0.16415683023634303   0.505620715124582   0.5468951671719203   0.6466441855491313   0.4644103619563068   0.6673279024590776   0.9205395790937742   0.7837633965476419
0.6481925280188677   0.471544798519523   0.16932271515606728   0.8893419605124154   0.30222073873881866   0.16485917971876393   0.5717462156842885   0.9786496400732295   0.6167464204968851   0.6036734846563317   0.1559262504231333   0.046402925046714096   0.22867957017185606   0.5264613715689335   0.8808204710863091   0.7441844116023881   0.06452273993551304   0.020840656444351534   0.3339253039143888   0.0975402260532568   0.6001123779792062   0.35351275398527393   0.41338572482061464   0.3137768295056148   0.9519198499603385   0.8819679554657509   0.2440630096645474   0.4244348689931994   0.6496991112215198   0.717108775746987   0.6723167939802589   0.44578522891996986   0.03295269072463472   0.11343529109065517   0.5163905435571257   0.39938230387325574   0.8042731205527787   0.5869739195217217   0.6355700724708164   0.6551978922708677   0.7397503806172656   0.5661332630773702   0.30164476855642763   0.5576576662176108   0.1396380026380594   0.2126205090920963   0.888259043735813   0.243880836711996   0.1877181526777209   0.3306525536263454   0.6441960340712656   0.8194459677187966   0.5380190414562012   0.6135437778793584   0.9718792400910067   0.3736607387988268   0.5050663507315664   0.5001084867887032   0.4554886965338811   0.9742784349255711   0.7007932301787877   0.9131345672669815   0.8199186240630646   0.3190805426547034
0.9610428495615221   0.3470013041896114   0.518273855506637   0.7614228764370926   0.8214048469234627   0.1343807950975151   0.630014811770824   0.5175420397250966   0.6336866942457418   0.8037282414711697   0.9858187776995584   0.6980960720063   0.09566765278954069   0.19018446359181126   0.013939537608551652   0.3244353332074732   0.5906013020579743   0.690075976803108   0.5584508410746706   0.35015689828190216   0.8898080718791865   0.7769414095361264   0.7385322170116059   0.031076355627198744   0.9287652223176645   0.42994010534651506   0.22025836150496894   0.2696534791901061   0.10736037539420175   0.29555931024899995   0.590243549734145   0.7521114394650096   0.4736736811484599   0.4918310687778303   0.6044247720345866   0.0540153674587096   0.3780060283589193   0.301646605186019   0.590485234426035   0.7295800342512364   0.7874047263009449   0.611570628382911   0.032034393351364376   0.37942313596933425   0.8975966544217584   0.8346292188467846   0.29350217633975845   0.3483467803421355   0.968831432104094   0.40468911350026954   0.07324381483478953   0.07869330115202934   0.8614710567098922   0.10912980325126954   0.4830002651006446   0.32658186168701975   0.38779737556143223   0.6172987344734393   0.878575493066058   0.27256649422831014   0.009791347202513   0.31565212928742026   0.2880902586400231   0.5429864599770737
0.22238662090156805   0.7040815009045093   0.2560558652886587   0.1635633240077395   0.3247899664798096   0.8694522820577246   0.9625536889489003   0.815216543665604   0.3559585343757157   0.4647631685574551   0.8893098741141107   0.7365232425135747   0.4944874776658235   0.35563336530618556   0.40630960901346613   0.4099413808265549   0.10669010210439124   0.7383346308327463   0.5277341159474082   0.13737488659824473   0.09689875490187824   0.42268250154532605   0.23964385730738505   0.594388426621171   0.8745121340003102   0.7186010006408168   0.9835879920187264   0.43082510261343143   0.5497221675205005   0.8491487185830922   0.021034303069826142   0.6156085589478274   0.19376363314478487   0.38438555002563707   0.13172442895571543   0.8790853164342527   0.6992761554789614   0.028752184719451478   0.7254148199422493   0.46914393560769785   0.5925860533745702   0.2904175538867052   0.1976807039948412   0.3317690490094531   0.4956872984726919   0.8677350523413792   0.9580368466874561   0.7373806223882821   0.6211751644723816   0.14913405170056238   0.9744488546687298   0.3065555197748506   0.07145299695188112   0.2999853331174702   0.9534145515989036   0.6909469608270232   0.8776893638070963   0.9155997830918332   0.8216901226431882   0.8118616443927705   0.17841320832813487   0.8868475983723817   0.09627530270093886   0.3427177087850727
0.5858271549535647   0.5964300444856765   0.8985945987060977   0.01094865977561958   0.09013985648087286   0.7286949921442973   0.9405577520186416   0.2735680373873375   0.46896469200849117   0.579560940443735   0.9661088973499118   0.9670125176124869   0.39751169505661005   0.27957560732626474   0.012694345751008189   0.2760655567854636   0.5198223312495138   0.3639758242344316   0.19100422310782   0.4642039123926931   0.3414091229213789   0.4771282258620499   0.09472892040688116   0.12148620360762045   0.7555819679678142   0.8806981813763733   0.1961343217007835   0.11053754383200087   0.6654421114869413   0.15200318923207606   0.25557656968214193   0.8369695064446634   0.19647741947845015   0.572442248788341   0.28946767233223014   0.8699569888321765   0.7989657244218401   0.2928666414620763   0.27677332658122195   0.593891432046713   0.27914339317232634   0.9288908172276448   0.08576910347340194   0.12968751965401987   0.9377342702509474   0.4517625913655948   0.9910401830665208   0.008201316046399402   0.18215230228313326   0.5710644099892215   0.7949058613657373   0.8976637722143985   0.516710190796192   0.4190612207571454   0.5393292916835953   0.060694265769735134   0.3202327713177418   0.8466189719688043   0.24986161935136522   0.19073727693755857   0.5212670468959016   0.553752330506728   0.9730882927701433   0.5968458448908456
0.2421236537235754   0.6248615132790832   0.8873191892967414   0.46715832523682577   0.30438938347262795   0.1730989219134884   0.8962790062302205   0.45895700919042637   0.12223708118949472   0.6020345119242669   0.10137314486448326   0.5612932369760278   0.6055268903933028   0.18297329116712155   0.5620438531808879   0.5005989712062927   0.285294119075561   0.3363543191983172   0.3121822338295227   0.3098616942687341   0.7640270721796593   0.7826019886915893   0.3390939410593794   0.7130158493778885   0.5219034184560839   0.15774047541250596   0.4517747517626381   0.24585752414106277   0.21751403498345595   0.9846415534990176   0.5554957455324175   0.7869005149506364   0.09527695379396121   0.3826070415747506   0.4541226006679343   0.22560727797460858   0.4897500634006584   0.1996337504076291   0.8920787474870464   0.725008306768316   0.20445594432509745   0.8632794312093118   0.5798965136575237   0.4151466124995818   0.44042887214543813   0.08067744251772266   0.24080257259814428   0.7021307631216933   0.9185254536893542   0.9229369671052167   0.7890278208355062   0.45627323898063055   0.7010114187058983   0.9382954136061991   0.23353207530308862   0.6693727240299941   0.605734464911937   0.5556883720314485   0.7794094746351543   0.44376544605538554   0.11598440151127866   0.3560546216238194   0.8873307271481079   0.7187571392870696
0.9115284571861813   0.4927751904145075   0.3074342134905842   0.3036105267874878   0.47109958504074306   0.4120977478967849   0.06663164089243993   0.6014797636657945   0.5525741313513888   0.48916078079156816   0.27760382005693374   0.14520652468516398   0.8515627126454905   0.550865367185369   0.04407174475384513   0.47583380065516984   0.24582824773355344   0.9951769951539206   0.2646622701186908   0.03206835459978433   0.12984384622227477   0.6391223735301012   0.37733154297058286   0.3133112153127147   0.21831538903609357   0.14634718311559367   0.06989732947999865   0.009700688525226897   0.7472158039953505   0.7342494352188088   0.00326568858755871   0.4082209248594324   0.19464167264396165   0.24508865442724065   0.725661868530625   0.2630144001742684   0.34307895999847116   0.6942232872418715   0.6815901237767799   0.7871805995190986   0.09725071226491769   0.699046292087951   0.41692785365808904   0.7551122449193143   0.9674068660426429   0.059923918557849815   0.039596310687506145   0.4418010296065995   0.7490914770065493   0.9135767354422561   0.9696989812075075   0.43210034108137263   0.0018756730111988622   0.1793273002234473   0.9664332926199488   0.023879416221940238   0.8072340003672372   0.9342386457962066   0.24077142408932384   0.7608650160476719   0.4641550403687661   0.2400153585543351   0.559181300312544   0.9736844165285733
0.3669043281038484   0.5409690664663841   0.142253446654455   0.21857217160925907   0.39949746206120545   0.48104514790853425   0.10265713596694885   0.7767711420026595   0.6504059850546561   0.5674684124662781   0.13295815475944137   0.34467080092128694   0.6485303120434572   0.3881411122428308   0.16652486213949258   0.3207913846993467   0.8412963116762201   0.45390246644662413   0.9257534380501687   0.5599263686516749   0.37714127130745395   0.21388710789228907   0.3665721377376247   0.5862419521231016   0.010236943203605603   0.672918041425905   0.22431869108316974   0.3676697805138425   0.6107394811424002   0.19187289351737072   0.12166155511622087   0.590898638511183   0.960333496087744   0.6244044810510926   0.9887034003567795   0.24622783758989603   0.3118031840442868   0.23626336880826176   0.8221785382172869   0.9254364528905493   0.47050687236806676   0.7823609023616376   0.8964251001671182   0.3655100842388745   0.09336560106061277   0.5684737944693485   0.5298529624294935   0.779268132115773   0.08312865785700717   0.8955557530434436   0.30553427134632377   0.4115983516019304   0.472389176714607   0.7036828595260729   0.1838727162301029   0.8206997130907475   0.512055680626863   0.07927837847498029   0.19516931587332337   0.5744718755008514   0.2002524965825762   0.8430150096667185   0.37299077765603644   0.6490354226103021
0.7297456242145095   0.060654107305080925   0.4765656774889182   0.28352533837142757   0.6363800231538966   0.4921803128357324   0.9467127150594247   0.5042572062556546   0.5532513652968896   0.5966245597922888   0.641178443713101   0.0926588546537242   0.08086218858228249   0.892941700266216   0.457305727482998   0.27195914156297674   0.5688065079554195   0.8136633217912357   0.26213641160967466   0.6974872660621253   0.36855401137284327   0.9706483121245172   0.8891456339536382   0.048451843451823184   0.6388083871583339   0.9099942048194363   0.41257995646472   0.7649265050803956   0.0024283640044371587   0.41781389198370383   0.4658672414052953   0.260669298824741   0.4491769987075476   0.821189332191415   0.8246887976921944   0.1680104441710168   0.3683148101252652   0.9282476319251991   0.3673830702091963   0.8960513026080401   0.7995083021698457   0.1145843101339634   0.10524665859952162   0.19856403654591478   0.43095429079700237   0.14393599800944626   0.21610102464588338   0.1501121930940916   0.7921459036386685   0.23394179319001004   0.8035210681811633   0.385185688013696   0.7897175396342314   0.8161279012063062   0.3376538267758681   0.12451638918895502   0.34054054092668373   0.9949385690148912   0.5129650290836737   0.9565059450179383   0.9722257308014186   0.06669093708969212   0.14558195887447742   0.060454642409898174
0.17271742863157288   0.9521066269557287   0.04033530027495581   0.8618906058639834   0.7417631378345705   0.8081706289462824   0.8242342756290725   0.7117784127698917   0.9496172341959019   0.5742288357562724   0.020713207447909075   0.3265927247561958   0.1598996945616706   0.7581009345499662   0.683059380672041   0.20207633556724075   0.8193591536349869   0.763162365535075   0.1700943515883673   0.24557039054930252   0.8471334228335683   0.6964714284453829   0.02451239271388986   0.18511574813940435   0.6744159942019954   0.7443648014896542   0.984177092438934   0.323225142275421   0.9326528563674249   0.9361941725433717   0.1599428168098616   0.6114467295055291   0.9830356221715228   0.3619653367870993   0.13922960936195253   0.28485400474933337   0.8231359276098523   0.6038644022371331   0.4561702286899115   0.08277766918209263   0.003776773974865445   0.8407020367020581   0.28607587710154425   0.8372072786327901   0.15664335114129715   0.14423060825667516   0.26156348438765437   0.6520915304933858   0.48222735693930174   0.399865806767021   0.27738639194872033   0.3288663882179648   0.5495745005718768   0.46367163422364926   0.11744357513885871   0.7174196587124356   0.566538878400354   0.10170629743654996   0.9782139657769062   0.43256565396310226   0.7434029507905017   0.49784189519941685   0.5220437370869947   0.3497879847810096
0.7396261768156362   0.6571398584973588   0.23596785998545042   0.5125807061482195   0.5829828256743391   0.5129092502406836   0.974404375597796   0.8604891756548337   0.10075546873503731   0.11304344347366262   0.6970179836490757   0.531622787436869   0.5511809681631604   0.6493718092500134   0.579574408510217   0.8142031287244333   0.9846420897628064   0.5476655118134633   0.6013604427333108   0.3816374747613311   0.24123913897230478   0.04982361661404653   0.07931670564631618   0.031849489980321465   0.5016129621566685   0.39268375811668776   0.8433488456608658   0.519268783832102   0.9186301364823295   0.8797745078760041   0.8689444700630697   0.6587796081772682   0.8178746677472921   0.7667310644023415   0.171926486413994   0.1271568207403993   0.26669369958413175   0.11735925515232817   0.592352077903777   0.312953692015966   0.28205160982132527   0.5696937433388648   0.9909916351704662   0.931316217254635   0.040812470849020496   0.5198701267248182   0.91167492952415   0.8994667272743134   0.5391995086923519   0.1271863686081305   0.06832608386328423   0.38019794344221153   0.6205693722100225   0.24741186073212637   0.19938161380021452   0.7214183352649433   0.8026947044627303   0.48068079632978483   0.02745512738622051   0.594261514524544   0.5360010048785986   0.3633215411774567   0.4351030494824435   0.28130782250857794
0.25394939505727326   0.7936277978385919   0.44411141431197737   0.349991605253943   0.21313692420825278   0.27375767111377364   0.5324364847878273   0.45052487797962953   0.6739374155159008   0.14657130250564315   0.46411040092454314   0.070326934537418   0.053368043305878396   0.8991594417735168   0.2647287871243286   0.34890859927247475   0.25067333884314813   0.4184786454437319   0.23727365973810813   0.7546470847479307   0.7146723339645495   0.05515710426627523   0.8021706102556646   0.47333926223935285   0.4607229389072763   0.26152930642768335   0.35805919594368724   0.12334765698540984   0.24758601469902347   0.9877716353139097   0.82562271115586   0.6728227790057804   0.5736485991831226   0.8412003328082666   0.36151231023131675   0.6024958444683624   0.5202805558772442   0.9420408910347497   0.09678352310698812   0.2535872451958876   0.2696072170340961   0.5235622455910178   0.85950986336888   0.4989401604479568   0.5549348830695465   0.46840514132474265   0.0573392531132154   0.025600898208603992   0.09421194416227031   0.2068758348970593   0.6992800571695281   0.9022532412231942   0.8466259294632468   0.21910419958314964   0.8736573460136683   0.2294304622174138   0.2729773302801242   0.3779038667748831   0.5121450357823515   0.6269346177490515   0.75269677440288   0.43586297574013333   0.41536151267536336   0.37334737255316386
0.48308955736878384   0.9123007301491155   0.5558516493064833   0.8744072121052071   0.9281546742992373   0.44389558882437286   0.4985123961932679   0.8488063138966031   0.833942730136967   0.23701975392731356   0.7992323390237398   0.9465530726734089   0.9873168006737201   0.017915554344163934   0.9255749930100715   0.7171226104559951   0.7143394703935959   0.6400116875692808   0.4134299572277201   0.09018799270694361   0.961642695990716   0.2041487118291475   0.9980684445523567   0.7168406201537797   0.4785531386219321   0.291847981680032   0.4422167952458734   0.8424334080485727   0.5503984643226949   0.8479523928556592   0.9437043990526054   0.9936270941519696   0.7164557341857279   0.6109326389283456   0.1444720600288656   0.047074021478560685   0.7291389335120078   0.5930170845841817   0.21889706701879402   0.3299514110225656   0.01479946311841188   0.9530053970149008   0.8054671097910739   0.23976341831562198   0.05315676712769592   0.7488566851857533   0.8073986652387173   0.5229227981618423   0.5746036285057637   0.4570087035057213   0.3651818699928439   0.6804893901132696   0.024205164183068926   0.6090563106500622   0.4214774709402385   0.6868622959613   0.307749429997341   0.9981236717217166   0.27700541091137293   0.6397882744827393   0.5786104964853332   0.4051065871375349   0.05810834389257889   0.3098368634601737
0.5638110333669213   0.4521011901226341   0.2526412341015049   0.07007344514455173   0.5106542662392254   0.7032445049368807   0.4452425688627877   0.5471506469827094   0.9360506377334616   0.24623580143115947   0.08006069886994374   0.8666612568694398   0.9118454735503927   0.6371794907810973   0.6585832279297053   0.1797989609081399   0.6040960435530517   0.6390558190593807   0.3815778170183323   0.5400106864254006   0.02548554706771847   0.23394923192184583   0.3234694731257534   0.2301738229652269   0.46167451370079715   0.7818480417992117   0.07082823902424848   0.16010037782067515   0.9510202474615718   0.07860353686233094   0.6255856701614608   0.6129497308379657   0.014969609728110126   0.8323677354311715   0.5455249712915171   0.7462884739685258   0.10312413617771744   0.19518824465007417   0.8869417433618119   0.5664895130603859   0.49902809262466574   0.5561324255906934   0.5053639263434795   0.026478826634985266   0.4735425455569473   0.3221831936688476   0.18189445321772613   0.7963050036697584   0.011868031856150152   0.5403351518696359   0.11106621419347765   0.6362046258490832   0.060847784394578414   0.4617316150073049   0.48548054403201685   0.023254895011117563   0.045878174666468284   0.6293638795761335   0.9399555727404998   0.2769664210425918   0.9427540384887508   0.43417563492605926   0.05301382937868793   0.7104769079822059
0.4437259458640851   0.8780432093353658   0.5476499030352084   0.6839980813472206   0.9701834003071378   0.5558600156665182   0.36575544981748226   0.8876930776774623   0.9583153684509876   0.015524863796882359   0.2546892356240046   0.25148845182837903   0.8974675840564093   0.5537932487895775   0.7692086915919878   0.22823355681726148   0.8515894093899409   0.924429369213444   0.829253118851488   0.9512671357746697   0.90883537090119   0.4902537342873847   0.7762392894728001   0.24079022779246378   0.465109425037105   0.6122105249520189   0.22858938643759172   0.5567921464452431   0.4949260247299672   0.05635050928550063   0.8628339366201094   0.6690990687677808   0.5366106562789796   0.04082564548861827   0.6081447009961048   0.4176106169394018   0.6391430722225704   0.48703239669904086   0.8389360094041171   0.18937706012214034   0.7875536628326294   0.5626030274855969   0.009682890552629036   0.23810992434747064   0.8787182919314394   0.07234929319821214   0.23344360107982895   0.9973196965550069   0.41360886689433435   0.46013876824619326   0.004854214642237235   0.44052755010976374   0.9186828421643671   0.40378825896069265   0.1420202780221278   0.7714284813419829   0.38207218588538755   0.36296261347207437   0.533875577026023   0.35381786440258106   0.7429291136628171   0.8759302167730335   0.6949395676219059   0.16444080428044075
0.9553754508301877   0.3133271892874367   0.6852566770692768   0.9263308799329701   0.07665715889874834   0.24097789608922454   0.4518130759894479   0.9290111833779633   0.663048292004414   0.7808391278430312   0.4469588613472107   0.4884836332681995   0.7443654498400468   0.37705086888233863   0.3049385833250829   0.7170551519262166   0.36229326395465933   0.014088255410264256   0.77106300629906   0.36323728752363554   0.6193641502918422   0.13815803863723072   0.07612343867715404   0.1987964832431948   0.6639886994616545   0.824830849349794   0.3908667616078772   0.2724656033102247   0.5873315405629062   0.5838529532605695   0.9390536856184293   0.34345441993226145   0.9242832485584921   0.8030138254175382   0.4920948242712186   0.854970786664062   0.17991779871844527   0.4259629565351996   0.18715624094613567   0.13791563473784535   0.8176245347637859   0.41187470112493535   0.4160932346470757   0.7746783472142098   0.19826038447194377   0.2737166624877046   0.33996979596992166   0.575881863971015   0.5342716850102893   0.4488858131379106   0.9491030343620445   0.30341626066079036   0.9469401444473832   0.8650328598773411   0.01004934874361524   0.9599618407285289   0.02265689588889106   0.06201903445980286   0.5179545244723966   0.10499105406446693   0.8427390971704458   0.6360560779246033   0.330798283526261   0.9670754193266216
0.025114562406659834   0.22418137679966793   0.9147050488791852   0.19239707211241175   0.826854177934716   0.9504647143119633   0.5747352529092636   0.6165152081413967   0.29258249292442673   0.5015789011740528   0.6256322185472191   0.3130989474806064   0.34564234847704356   0.6365460412967117   0.6155828698036039   0.3531371067520775   0.3229854525881525   0.5745270068369088   0.09762834533120718   0.24814605268761059   0.4802463554177067   0.9384709289123055   0.7668300618049462   0.28107063336098903   0.45513179301104684   0.7142895521126376   0.8521250129257609   0.08867356124857725   0.6282776150763308   0.7638248378006742   0.27738976001649734   0.4721583531071805   0.33569512215190406   0.26224593662662155   0.6517575414692782   0.1590594056265741   0.9900527736748606   0.6256998953299099   0.036174671665674396   0.8059222988744966   0.6670673210867081   0.051172888493001056   0.9385463263344672   0.557776246186886   0.18682096566900136   0.11270195958069554   0.17171626452952105   0.276705612825897   0.7316891726579545   0.39841240746805795   0.3195912516037601   0.18803205157731975   0.10341155758162368   0.6345875696673837   0.04220149158726279   0.7158736984701393   0.7677164354297196   0.3723416330407622   0.39044395011798455   0.5568142928435651   0.7776636617548591   0.7466417377108523   0.35426927845231015   0.7508919939690685
0.11059634066815105   0.6954688492178512   0.41572295211784294   0.19311574778218246   0.9237753749991497   0.5827668896371557   0.2440066875883219   0.9164101349562854   0.19208620234119522   0.18435448216909778   0.9244154359845618   0.7283780833789657   0.08867464475957153   0.5497669125017141   0.8822139443972989   0.012504384908826447   0.3209582093298519   0.17742527946095193   0.49176999427931445   0.45569009206526134   0.5432945475749928   0.43078354175009964   0.1375007158270043   0.7047980980961929   0.43269820690684174   0.7353146925322483   0.7217777637091614   0.5116823503140103   0.508922831907692   0.15254780289509268   0.47777107612083947   0.5952722153577249   0.31683662956649683   0.968193320725995   0.5533556401362777   0.8668941319787592   0.22816198480692532   0.41842640822428084   0.6711416957389786   0.8543897470699328   0.9072037754770734   0.2410011287633289   0.17937170145966425   0.3986996550046714   0.36390922790208063   0.8102175870132293   0.04187098563265996   0.6939015569084787   0.9312110209952389   0.07490289448098088   0.3200932219234986   0.18221920659446825   0.4222881890875468   0.9223550915858882   0.8423221458026592   0.5869469912367433   0.10545155952104997   0.9541617708598933   0.2889665056663815   0.7200528592579841   0.8772895747141246   0.5357353626356125   0.6178248099274027   0.8656631121880514
0.9700857992370512   0.2947342338722836   0.43845310846773855   0.4669634571833799   0.6061765713349706   0.4845166468590543   0.3965821228350786   0.7730619002749013   0.6749655503397317   0.4096137523780734   0.07648890091157998   0.5908426936804331   0.25267736125218493   0.4872586607921852   0.23416675510892082   0.003895702443689711   0.14722580173113498   0.5330968899322919   0.9452002494425393   0.2838428431857056   0.2699362270170103   0.9973615272966795   0.32737543951513653   0.4181797309976542   0.29985042777995913   0.7026272934243959   0.888922331047398   0.9512162738142743   0.6936738564449885   0.21811064656534157   0.49234020821231944   0.17815437353937302   0.01870830610525677   0.8084968941872681   0.41585130730073944   0.58731167985894   0.7660309448530719   0.3212382333950829   0.18168455219181864   0.5834159774152503   0.6188051431219369   0.788141343462791   0.23648430274927928   0.2995731342295447   0.34886891610492654   0.7907798161661116   0.9091088632341428   0.8813934032318904   0.04901848832496741   0.08815252274171567   0.02018653218674471   0.9301771294176161   0.3553446318799789   0.8700418761763741   0.5278463239744253   0.7520227558782431   0.33663632577472213   0.06154498198910599   0.11199501667368582   0.16471107601930313   0.5706053809216503   0.7403067485940231   0.9303104644818672   0.5812950986040528
0.9518002377997135   0.952165405131232   0.6938261617325879   0.2817219643745082   0.6029313216947869   0.16138558896512054   0.7847172984984452   0.4003285611426178   0.5539128333698194   0.07323306622340486   0.7645307663117005   0.4701514317250017   0.19856820148984058   0.20319119004703073   0.23668444233727517   0.7181286758467585   0.8619318757151184   0.14164620805792477   0.12468942566358936   0.5534175998274554   0.29132649479346817   0.4013394594639017   0.19437896118172218   0.9721225012234026   0.3395262569937547   0.4491740543326696   0.5005527994491343   0.6904005368488944   0.7365949352989678   0.28778846536754904   0.7158355009506892   0.2900719757062766   0.1826821019291483   0.2145553991441442   0.9513047346389887   0.8199205439812749   0.9841139004393077   0.011364209097113446   0.7146202923017135   0.10179186813451639   0.12218202472418926   0.8697180010391887   0.5899308666381242   0.5483742683070609   0.8308555299307211   0.468378541575287   0.395551905456402   0.5762517670836584   0.49132927293696643   0.0192044872426174   0.8949991060072677   0.8858512302347641   0.7547343376379986   0.7314160218750684   0.17916360505657855   0.5957792545284875   0.5720522357088503   0.5168606227309241   0.22785887041758984   0.7758587105472124   0.5879383352695426   0.5054964136338107   0.5132385781158764   0.6740668424126961
0.4657563105453533   0.635778412594622   0.9233077114777521   0.12569257410563514   0.6349007806146323   0.167399871019335   0.5277558060213502   0.5494408070219767   0.14357150767766583   0.14819538377671762   0.6327567000140825   0.6635895767872128   0.3888371700396672   0.41677936190164927   0.45359309495750394   0.06781032225872528   0.8167849343308169   0.8999187391707252   0.2257342245399141   0.2919516117115128   0.2288465990612743   0.3944223255369144   0.7124956464240378   0.6178847692988166   0.763090288515921   0.7586439129422924   0.7891879349462857   0.4921921951931815   0.12818950790128872   0.5912440419229574   0.2614321289249355   0.9427513881712049   0.9846180002236229   0.4430486581462398   0.628675428910853   0.2791618113839921   0.5957808301839557   0.026269296244590505   0.17508233395334905   0.2113514891252668   0.7789958958531388   0.1263505570738654   0.949348109413435   0.9193998774137541   0.5501492967918644   0.731928231536951   0.23685246298939716   0.3015151081149373   0.7870590082759436   0.9732843185946586   0.4476645280431115   0.8093229129217557   0.6588695003746547   0.38204027667170115   0.18623239911817605   0.866571524750551   0.674251500151032   0.9389916185254613   0.5575569702073231   0.5874097133665589   0.07847066996707626   0.9127223222808709   0.382474636253974   0.3760582242412921
0.29947477411393747   0.7863717652070055   0.43312652684053904   0.45665834682753803   0.749325477322073   0.05444353367005453   0.19627406385114188   0.15514323871260072   0.9622664690461296   0.08115921507539599   0.7486095358080304   0.34582032579084493   0.30339696867147475   0.6991189384036949   0.5623771366898543   0.47924880104029394   0.6291454685204428   0.7601273198782335   0.004820166482531279   0.8918390876737351   0.5506747985533665   0.8474049975973627   0.6223455302285573   0.515780863432443   0.25120002443942907   0.06103323239035713   0.18921900338801828   0.05912251660490494   0.501874547117356   0.0065896987203025986   0.9929449395368763   0.9039792778923043   0.5396080780712265   0.9254304836449067   0.24433540372884605   0.5581589521014593   0.23621110939975176   0.22631154524121178   0.6819582670389918   0.07891015106116532   0.6070656408793089   0.4661842253629783   0.6771381005564605   0.18707106338743026   0.056390842325942395   0.6187792277656157   0.05479257032790316   0.6712901999549873   0.8051908178865134   0.5577459953752586   0.8655735669398849   0.6121676833500823   0.3033162707691573   0.551156296654956   0.8726286274030085   0.7081884054577782   0.7637081926979308   0.6257258130100494   0.6282932236741624   0.15002945335631884   0.527497083298179   0.3994142677688376   0.9463349566351708   0.07111930229515351
0.9204314424188701   0.9332300424058593   0.26919685607871024   0.8840482389077232   0.8640406000929277   0.31445081464024355   0.21440428575080708   0.21275803895273598   0.05884978220641433   0.756704819264985   0.3488307188109222   0.6005903556026536   0.755533511437257   0.20554852261002898   0.4762020914079137   0.8924019501448756   0.9918253187393262   0.5798227095999796   0.8479088677337513   0.7423724967885567   0.4643282354411472   0.18040844183114202   0.9015739110985805   0.6712531944934031   0.5438967930222771   0.24717839942528275   0.6323770550198703   0.7872049555856799   0.6798561929293495   0.9327275847850391   0.41797276926906324   0.574446916632944   0.6210064107229352   0.17602276552005422   0.06914205045814105   0.9738565610302903   0.8654728992856782   0.9704742429100253   0.5929399590502273   0.0814546108854148   0.8736475805463519   0.39065153331004565   0.745031091316476   0.3390821140968581   0.4093193451052047   0.2102430914789036   0.8434571802178955   0.6678289196034549   0.8654225520829275   0.9630646920536209   0.21108012519802516   0.880623964017775   0.18556635915357803   0.030337107268581655   0.7931073559289619   0.30617704738483104   0.5645599484306428   0.8543143417485274   0.7239653054708208   0.3323204863545407   0.6990870491449648   0.8838400988385022   0.13102534642059352   0.2508658754691259
0.8254394685986128   0.4931885655284566   0.38599425510411745   0.9117837613722678   0.41612012349340816   0.28294547404955295   0.5425370748862219   0.24395484176881288   0.5506975714104807   0.3198807819959321   0.3314569496881968   0.3633308777510379   0.36513121225690265   0.2895436747273505   0.5383495937592349   0.05715383036620685   0.8005712638262598   0.43522933297882305   0.814384288288414   0.7248333440116661   0.10148421468129501   0.5513892341403208   0.6833589418678205   0.47396746854254024   0.27604474608268215   0.05820066861186427   0.29736468676370303   0.5621837071702724   0.8599246225892739   0.7752551945623113   0.754827611877481   0.31822886540145956   0.3092270511787933   0.45537441256637917   0.42337066218928426   0.9548979876504217   0.9440958389218906   0.16583073783902874   0.8850210684300495   0.8977441572842149   0.14352457509563094   0.7306014048602057   0.0706367801416354   0.17291081327254867   0.04204036041433592   0.17921217071988488   0.3872778382738149   0.6989433447300084   0.7659956143316538   0.1210115021080206   0.08991315151011187   0.13675963755973602   0.9060709917423798   0.3457563075457093   0.33508553963263077   0.8185307721582765   0.5968439405635865   0.8903818949793301   0.9117148774433464   0.8636327845078549   0.6527481016416958   0.7245511571403014   0.02669380901329708   0.96588862722364
0.5092235265460648   0.9939497522800956   0.9560570288716617   0.7929778139510913   0.46718316613172894   0.8147375815602108   0.5687791905978468   0.0940344692210829   0.7011875518000752   0.6937260794521902   0.47886603908773495   0.9572748316613469   0.7951165600576954   0.3479697719064809   0.14378049945510415   0.1387440595030704   0.1982726194941089   0.4575878769271508   0.23206562201175765   0.27511127499521554   0.5455245178524131   0.7330367197868495   0.20537181299846058   0.30922264777157554   0.03630099130634822   0.7390869675067537   0.2493147841267989   0.5162448338204841   0.5691178251746193   0.924349385946543   0.6805355935289521   0.4222103645994013   0.8679302733745441   0.2306233064943528   0.20166955444121717   0.4649355329380544   0.07281371331684872   0.8826535345878719   0.05788905498611303   0.326191473434984   0.8745410938227398   0.42506565766072113   0.8258234329743553   0.051080198439768465   0.32901657597032674   0.6920289378738718   0.6204516199758948   0.7418575506681929   0.2927155846639785   0.9529419703671179   0.3711368358490959   0.22561271684770873   0.7235977594893592   0.028592584420574947   0.6906012423201437   0.8034023522483075   0.8556674861148151   0.7979692779262222   0.4889316878789266   0.338466819310253   0.7828537727979664   0.9153157433383502   0.4310426328928136   0.012275345875269014
0.9083126789752266   0.49025008567762907   0.6052191999184582   0.9611951474355005   0.5792961030048999   0.7982211478037573   0.9847675799425635   0.21933759676730763   0.2865805183409214   0.8452791774366394   0.6136307440934675   0.9937248799195989   0.5629827588515621   0.8166865930160645   0.9230295017733238   0.19032252767129143   0.7073152727367471   0.018717315089842316   0.43409781389439717   0.8518557083610384   0.9244614999387807   0.10340157175149212   0.0030551810015835784   0.8395803624857694   0.01614882096355405   0.613151486073863   0.39783598108312535   0.8783852150502688   0.43685271795865416   0.8149303382701057   0.4130684011405619   0.6590476182829612   0.15027219961773278   0.9696511608334664   0.7994376570470945   0.6653227383633623   0.5872894407661706   0.15296456781740186   0.8764081552737707   0.4750002106920709   0.8799741680294235   0.13424725272755955   0.44231034137937353   0.6231445023310325   0.9555126680906428   0.030845680976067436   0.43925516037778994   0.7835641398452631   0.9393638471270889   0.4176941949022044   0.04141917929466455   0.9051789247949943   0.5025111291684347   0.6027638566320986   0.6283507781541026   0.24613130651203305   0.3522389295507019   0.6331126957986324   0.8289131211070082   0.5808085681486708   0.7649494887845313   0.48014812798123047   0.9525049658332375   0.10580835745659985
0.8849753207551078   0.3459008752536709   0.5101946244538641   0.48266385512556736   0.9294626526644649   0.3150551942776035   0.07093946407607413   0.6990997152803042   0.9900988055373761   0.8973609993753991   0.02952028478140957   0.79392079048531   0.4875876763689414   0.29459714274330046   0.40116950662730694   0.547789483973277   0.1353487468182395   0.6614844469446681   0.5722563855202988   0.9669809158246062   0.37039925803370816   0.18133631896343763   0.6197514196870613   0.8611725583680064   0.4854239372786004   0.8354354437097667   0.10955679523319717   0.378508703242439   0.5559612846141355   0.5203802494321632   0.038617331157123055   0.6794089879621348   0.5658624790767595   0.6230192500567641   0.009097046375713482   0.8854881974768247   0.07827480270781807   0.32842210731346366   0.6079275397484065   0.3376987135035478   0.9429260558895786   0.6669376603687955   0.03567115422810776   0.3707177976789416   0.5725267978558705   0.48560134140535793   0.4159197345410465   0.5095452393109352   0.08710286057727   0.6501658976955913   0.30636293930784936   0.1310365360684962   0.5311415759631345   0.12978564826342803   0.2677456081507263   0.4516275481063614   0.965279096886375   0.5067663982066639   0.25864856177501283   0.5661393506295367   0.887004294178557   0.17834429089320028   0.6507210220266063   0.22844063712598883
0.9440782382889784   0.5114066305244047   0.6150498677984986   0.8577228394470472   0.37155144043310795   0.025805289119046795   0.19913013325745202   0.34817760013611204   0.28444857985583794   0.37563939142345554   0.8927671939496027   0.21714106406761582   0.7533070038927034   0.2458537431600275   0.6250215857988763   0.7655135159612544   0.7880279070063284   0.7390873449533636   0.3663730240238635   0.19937416533171773   0.9010236128277714   0.5607430540601632   0.7156520019972572   0.9709335282057289   0.9569453745387931   0.04933642353575853   0.10060213419875866   0.11321068875868165   0.5853939341056852   0.023531134416711733   0.9014720009413066   0.7650330886225696   0.30094535424984725   0.6478917429932561   0.008704806991703985   0.5478920245549538   0.5476383503571438   0.4020379998332287   0.38368322119282766   0.7823785085936994   0.7596104433508153   0.6629506548798652   0.017310197168964127   0.5830043432619817   0.8585868305230439   0.10220760081970186   0.30165819517170694   0.6120708150562528   0.9016414559842507   0.05287117728394333   0.20105606097294826   0.4988601262975711   0.3162475218785656   0.0293400428672316   0.2995840600316416   0.7338270376750015   0.01530216762871835   0.3814482998739754   0.29087925303993767   0.18593501312004768   0.4676638172715746   0.9794103000407467   0.90719603184711   0.4035565045263483
0.7080533739207593   0.3164596451608816   0.8898858346781459   0.8205521612643666   0.8494665433977153   0.21425204434117973   0.588227639506439   0.20848134620811384   0.9478250874134646   0.1613808670572364   0.3871715785334907   0.7096212199105427   0.6315775655348991   0.13204082419000482   0.08758751850184905   0.9757941822355413   0.6162753979061807   0.7505925243160294   0.7967082654619114   0.7898591691154936   0.1486115806346061   0.7711822242752827   0.8895122336148014   0.38630266458914525   0.4405582067138469   0.45472257911440106   0.9996263989366555   0.5657505033247786   0.5910916633161315   0.24047053477322133   0.4113987594302166   0.3572691571166648   0.6432665759026669   0.07908966771598493   0.024227180896725896   0.647647937206122   0.01168901036776784   0.9470488435259802   0.9366396623948768   0.6718537549705809   0.3954136124615871   0.1964563192099507   0.13993139693296544   0.8819945858550873   0.24680203182698102   0.42527409493466806   0.250419163318164   0.495691921265942   0.8062438251131341   0.970551515820267   0.2507927643815085   0.9299414179411634   0.21515216179700264   0.7300809810470457   0.8393940049512919   0.5726722608244986   0.5718855858943357   0.6509913133310608   0.815166824054566   0.9250243236183765   0.5601965755265679   0.7039424698050806   0.8785271616596891   0.2531705686477957
0.16478296306498075   0.5074861505951299   0.7385957647267237   0.3711759827927084   0.9179809312379997   0.08221205566046182   0.48817660140855973   0.8754840615267664   0.11173710612486559   0.11166053984019483   0.23738383702705124   0.9455426435856029   0.896584944327863   0.3815795587931492   0.39798983207575933   0.37287038276110435   0.3246993584335272   0.7305882454620884   0.5828230080211934   0.4478460591427278   0.7645027829069594   0.026645775657007858   0.7042958463615041   0.1946754904949321   0.5997198198419785   0.519159625061878   0.9657000816347804   0.8234995077022237   0.6817388886039788   0.43694756940141616   0.4775234802262207   0.9480154461754573   0.5700017824791133   0.32528702956122135   0.24013964319916944   0.0024728025898543725   0.6734168381512503   0.9437074707680722   0.8421498111234101   0.62960241982875   0.34871747971772304   0.2131192253059837   0.2593268031022168   0.18175636068602224   0.5842146968107637   0.18647344964897586   0.5550309567407126   0.9870808701910901   0.9844948769687851   0.6673138245870979   0.5893308751059322   0.16358136248886646   0.30275598836480627   0.23036625518568168   0.11180739487971153   0.21556591631340913   0.7327542058856931   0.9050792256244603   0.8716677516805421   0.21309311372355477   0.05933736773444276   0.9613717548563881   0.029517940557131972   0.5834906938948047
0.7106198880167197   0.7482525295504044   0.7701911374549152   0.4017343332087825   0.12640519120595603   0.5617790799014286   0.21516018071420256   0.41465346301769235   0.1419103142371709   0.8944652553143307   0.6258293056082703   0.2510721005288259   0.8391543258723646   0.6640990001286491   0.5140219107285589   0.03550618421541675   0.10640011998667158   0.7590197745041888   0.6423541590480167   0.822413070491862   0.047062752252228814   0.7976480196478005   0.6128362184908848   0.23892237659705726   0.33644286423550906   0.049395490097396064   0.8426450810359696   0.8371880433882748   0.21003767302955306   0.4876164101959674   0.6274849003217671   0.42253458037058245   0.06812735879238219   0.5931511548816366   0.0016555947134966516   0.17146247984175655   0.22897303292001758   0.9290521547529875   0.4876336839849378   0.1359562956263398   0.122572912933346   0.17003238024879885   0.845279524936921   0.3135432251344778   0.07551016068111718   0.3723843606009983   0.23244330644603625   0.07462084853742054   0.7390672964456081   0.32298887050360225   0.38979822541006665   0.23743280514914578   0.529029623416055   0.8353724603076348   0.7623133250882996   0.8148982247785633   0.46090226462367284   0.24222130542599812   0.760657730374803   0.6434357449368068   0.23192923170365526   0.31316915067301054   0.27302404638986516   0.507479449310467
0.10935631877030927   0.14313677042421172   0.4277445214529441   0.19393622417598919   0.033846158089192085   0.7707524098232135   0.1953012150069079   0.11931537563856864   0.29477886164358397   0.4477635393196112   0.8055029895968412   0.8818825704894229   0.7657492382275289   0.6123910790119764   0.04318966450854157   0.06698434571085954   0.30484697360385615   0.37016977358597825   0.28253193413373856   0.42354860077405276   0.07291774190020087   0.0570006229129677   0.009507887743873395   0.9160691514635858   0.9635614231298916   0.913863852488756   0.5817633662909293   0.7221329272875966   0.9297152650406995   0.14311144266554257   0.3864621512840214   0.602817551649028   0.6349364033971155   0.6953479033459313   0.5809591616871802   0.7209349811596051   0.8691871651695865   0.08295682433395496   0.5377694971786385   0.6539506354487455   0.5643401915657305   0.7127870507479767   0.2552375630449   0.23040203467469278   0.49142244966552956   0.655786427835009   0.2457296753010266   0.314332883211107   0.5278610265356379   0.741922575346253   0.6639663090100973   0.5921999559235104   0.5981457614949385   0.5988111326807104   0.27750415772607595   0.9893824042744824   0.9632093580978229   0.9034632293347791   0.6965449960388959   0.26844742311487735   0.09402219292823638   0.8205064050008242   0.15877549886025724   0.6144967876661318
0.529682001362506   0.10771935425284744   0.9035379358153572   0.384094752991439   0.03825955169697642   0.45193292641783844   0.6578082605143306   0.06976186978033205   0.5103985251613384   0.7100103510715854   0.9938419515042333   0.4775619138568217   0.9122527636664001   0.11119921839087497   0.7163377937781573   0.4881795095823392   0.9490434055685771   0.2077359890560959   0.019792797739261486   0.21973208646746187   0.8550212126403407   0.38722958405527175   0.8610172988790042   0.6052352988013301   0.3253392112778347   0.27951022980242435   0.957479363063647   0.22114054580989098   0.2870796595808583   0.8275773033845859   0.29967110254931634   0.15137867602955896   0.7766811344195198   0.11756695231300045   0.30582915104508307   0.6738167621727373   0.8644283707531198   0.006367733922125466   0.5894913572669257   0.18563725259039807   0.9153849651845427   0.7986317448660296   0.5696985595276642   0.9659051661229362   0.06036375254420205   0.4114021608107578   0.70868126064866   0.36066986732160616   0.7350245412663673   0.1318919310083335   0.751201897585013   0.13952932151171518   0.447944881685509   0.3043146276237476   0.45153079503569665   0.9881506454821563   0.6712637472659891   0.18674767531074718   0.1457016439906136   0.31433388330941897   0.8068353765128693   0.1803799413886217   0.5562102867236879   0.12869663071902088
0.8914504113283266   0.3817481965225921   0.9865117271960236   0.16279146459608465   0.8310866587841245   0.9703460357118343   0.2778304665473636   0.8021215972744785   0.09606211751775716   0.8384541047035008   0.5266285689623506   0.6625922757627632   0.6481172358322481   0.5341394770797532   0.07509777392665389   0.674441630280607   0.976853488566259   0.347391801769006   0.9293961299360403   0.3601077469711881   0.17001811205338974   0.16701186038038432   0.37318584321235243   0.2314111162521672   0.2785677007250632   0.7852636638577922   0.3866741160163288   0.06861965165608255   0.4474810419409387   0.8149176281459579   0.10884364946896521   0.26649805438160407   0.35141892442318157   0.976463523442457   0.5822150805066146   0.6039057786188408   0.7033016885909333   0.4423240463627039   0.5071173065799608   0.9294641483382338   0.7264482000246744   0.09493224459369784   0.5777211766439205   0.5693564013670457   0.5564300879712846   0.9279203842133136   0.2045353334315681   0.3379452851148784   0.2778623872462214   0.14265672035552135   0.8178612174152393   0.2693256334587959   0.8303813453052827   0.3277390922095635   0.7090175679462741   0.0028275790771918217   0.47896242088210117   0.3512755687671064   0.12680248743965944   0.398921800458351   0.7756607322911678   0.9089515224044026   0.6196851808596986   0.4694576521201173
0.049212532266493456   0.8140192778107047   0.04196400421577813   0.9001012507530717   0.49278244429520884   0.8860988935973911   0.83742867078421   0.5621559656381933   0.2149200570489874   0.7434421732418698   0.019567453368970703   0.2928303321793973   0.3845387117437047   0.41570308103230635   0.3105498854226966   0.29000275310220547   0.9055762908616035   0.06442751226519994   0.1837473979830372   0.8910809526438545   0.12991555857043569   0.1554759898607974   0.5640622171233385   0.42162330052373714   0.08070302630394223   0.3414567120500927   0.5220982129075604   0.5215220497706655   0.5879205820087334   0.4553578184527015   0.6846695421233504   0.9593660841324723   0.373000524959746   0.7119156452108317   0.6651020887543797   0.666535751953075   0.9884618132160413   0.2962125641785253   0.3545522033316831   0.3765329988508695   0.08288552235443782   0.2317850519133254   0.1708048053486459   0.48545204620701504   0.9529699637840021   0.076309062052528   0.6067425882253074   0.06382874568327787   0.8722669374800599   0.7348523500024353   0.08464437531774696   0.5423066959126124   0.28434635547132653   0.2794945315497338   0.3999748331943966   0.5829406117801401   0.9113458305115805   0.5675788863389021   0.7348727444400169   0.9164048598270651   0.9228840172955391   0.2713663221603768   0.3803205411083338   0.5398718609761957
0.8399984949411013   0.039581270247051395   0.2095157357596879   0.0544198147691806   0.8870285311570992   0.9632722081945234   0.6027731475343805   0.9905910690859028   0.014761593677039355   0.22841985819208804   0.5181287722166336   0.44828437317329034   0.7304152382057129   0.9489253266423543   0.118153939022237   0.8653437613931503   0.8190694076941324   0.3813464403034521   0.38328119458222015   0.9489389015660852   0.8961853903985931   0.10998011814307532   0.002960653473886324   0.4090670405898896   0.05618689545749177   0.07039884789602392   0.7934449177141984   0.35464722582070896   0.16915836430039252   0.10712663970150053   0.19067177017981787   0.36405615673480624   0.15439677062335316   0.8787067815094125   0.6725429979631843   0.9157717835615159   0.4239815324176403   0.9297814548670582   0.5543890589409473   0.05042802216836558   0.604912124723508   0.5484350145636061   0.17110786435872716   0.10148912060228041   0.7087267343249148   0.4384548964205308   0.16814721088484083   0.6924220800123908   0.6525398388674231   0.3680560485245069   0.3747022931706424   0.3377748541916819   0.4833814745670305   0.26092940882300636   0.18403052299082454   0.9737186974568757   0.32898470394367735   0.38222262731359385   0.5114875250276403   0.05794691389535984   0.905003171526037   0.45244117244653564   0.9570984660866929   0.007518891726994256
0.3000910468025291   0.9040061578829295   0.7859906017279658   0.9060297711247138   0.5913643124776142   0.46555126146239867   0.6178433908431249   0.213607691112323   0.9388244736101913   0.09749521293789179   0.24314109767248251   0.8758328369206411   0.4554429990431607   0.8365658041148855   0.059110574681657965   0.9021141394637654   0.12645829509948334   0.45434317680129155   0.5476230496540178   0.8441672255684055   0.22145512357344627   0.0019020043547559044   0.5905245835673247   0.8366483338414112   0.9213640767709171   0.09789584647182639   0.804533981839359   0.9306185627166974   0.32999976429330286   0.6323445850094277   0.18669059099623408   0.7170108716043745   0.39117529068311163   0.5348493720715359   0.9435494933237516   0.8411780346837334   0.935732291639951   0.6982835679566505   0.8844389186420936   0.939063895219968   0.8092739965404676   0.24394039115535895   0.33681586898807586   0.09489666965156245   0.5878188729670214   0.24203838680060305   0.7462912854207511   0.25824833581015116   0.6664547961961041   0.14414254032877666   0.9417573035813921   0.3276297730934537   0.3364550319028013   0.5117979553193489   0.755066712585158   0.6106189014890793   0.9452797412196896   0.976948583247813   0.8115172192614064   0.7694408668053458   0.009547449579738715   0.2786650152911625   0.9270783006193128   0.8303769715853779
0.2002734530392711   0.03472462413580356   0.5902624316312369   0.7354803019338154   0.6124545800722497   0.7926862373352005   0.8439711462104859   0.4772319661236643   0.9459997838761456   0.6485436970064239   0.9022138426290938   0.14960219303021058   0.6095447519733442   0.1367457416870749   0.1471471300439358   0.5389832915411313   0.6642650107536546   0.1597971584392619   0.33562991078252935   0.7695424247357854   0.6547175611739159   0.8811321431480994   0.40855161016321656   0.9391654531504074   0.4544441081346448   0.8464075190122958   0.8182891785319797   0.20368515121659203   0.841989528062395   0.05372128167709531   0.9743180323214938   0.7264531850929278   0.8959897441862494   0.40517758467067144   0.07210418969240004   0.5768509920627172   0.2864449922129052   0.26843184298359657   0.9249570596484643   0.03786770052158587   0.6221799814592506   0.10863468454433466   0.5893271488659348   0.26832527578580045   0.9674624202853347   0.22750254139623527   0.18077553870271834   0.32915982263539295   0.5130183121506899   0.38109502238393944   0.3624863601707387   0.12547467141880092   0.6710287840882948   0.32737374070684416   0.3881683278492449   0.3990214863258732   0.7750390399020454   0.9221961560361727   0.31606413815684486   0.822170494263156   0.48859404768914017   0.6537643130525761   0.3911070785083806   0.7843027937415702
0.8664140662298896   0.5451296285082414   0.8017799296424457   0.5159775179557696   0.8989516459445549   0.3176270871120062   0.6210043909397274   0.1868176953203767   0.385933333793865   0.9365320647280667   0.25851803076898866   0.061343023901575776   0.7149045497055702   0.6091583240212226   0.8703497029197438   0.6623215375757026   0.9398655098035248   0.6869621679850499   0.5542855647628989   0.8401510433125465   0.4512714621143846   0.033197854932473805   0.16317848625451833   0.05584824957097642   0.584857395884495   0.4880682264242323   0.36139855661207265   0.5398707316152067   0.6859057499399401   0.17044113931222615   0.7403941656723453   0.35305303629483004   0.29997241614607506   0.2339090745841594   0.4818761349033566   0.2917100123932543   0.5850678664405049   0.6247507505629368   0.6115264319836128   0.6293884748175517   0.6452023566369801   0.9377885825778869   0.05724086722071389   0.7892374315050051   0.19393089452259543   0.904590727645413   0.8940623809661955   0.7333891819340287   0.6090734986381005   0.41652250122118073   0.532663824354123   0.19351845031882195   0.9231677486981603   0.24608136190895458   0.7922696586817777   0.8404654140239919   0.6231953325520853   0.012172287324795176   0.31039352377842105   0.5487554016307377   0.038127466111580334   0.38742153676185836   0.6988670917948082   0.919366926813186
0.39292510947460024   0.44963295418397153   0.6416262245740944   0.13012949530818088   0.19899421495200484   0.5450422265385585   0.7475638436078987   0.39674031337415216   0.5899207163139044   0.12851972531737774   0.21490001925377586   0.20322186305533024   0.6667529676157441   0.8824383634084232   0.4226303605719982   0.36275644903133836   0.04355763506365892   0.870266076083628   0.11223683679357718   0.8140010474006008   0.005430168952078586   0.48284453932176963   0.413369744998769   0.8946341205874148   0.6125050594774784   0.033211585137798094   0.7717435204246746   0.7645046252792339   0.4135108445254735   0.48816935859923966   0.024179676816775894   0.3677643119050817   0.8235901282115691   0.3596496332818619   0.809279657563   0.16454244884975142   0.15683716059582492   0.4772112698734387   0.3866492969910018   0.801785999818413   0.11327952553216601   0.6069451937898107   0.27441246019742466   0.9877849524178124   0.10784935658008742   0.1241006544680411   0.8610427151986557   0.09315083183039764   0.4953442971026091   0.090889069330243   0.089299194773981   0.3286462065511638   0.0818334525771356   0.6027197107310034   0.06511951795720511   0.9608818946460821   0.2582433243655666   0.2430700774491415   0.2558398603942051   0.7963394457963308   0.10140616376974163   0.7658588075757028   0.8691905634032032   0.9945534459779176
0.9881266382375756   0.15891361378589205   0.5947781032057786   0.006768493560105276   0.8802772816574882   0.03481295931785096   0.7337353880071229   0.9136176617297076   0.3849329845548791   0.9439238899876079   0.6444361932331419   0.5849714551785439   0.3030995319777435   0.34120417925660457   0.5793166752759368   0.6240895605324617   0.044856207612176936   0.09813410180746308   0.32347681488173174   0.827750114736131   0.9434500438424354   0.3322752942317603   0.4542862514785285   0.8331966687582133   0.9553234056048597   0.17336168044586822   0.8595081482727499   0.8264281751981081   0.0750461239473715   0.13854872112801728   0.12577276026562698   0.9128105134684005   0.6901131393924924   0.19462483114040932   0.48133656703248506   0.3278390582898566   0.38701360741474894   0.8534206518838048   0.9020198917565482   0.7037494977573949   0.342157399802572   0.7552865500763417   0.5785430768748164   0.8759993830212639   0.3987073559601367   0.4230112558445814   0.12425682539628793   0.042802714263050545   0.44338395035527695   0.24964957539871313   0.264748677123538   0.21637453906494247   0.36833782640790547   0.11110085427069587   0.13897591685791102   0.30356402559654205   0.678224687015413   0.9164760231302865   0.657639349825426   0.9757249673066855   0.2912110796006641   0.0630553712464818   0.7556194580688778   0.2719754695492905
0.9490536797980922   0.30776882117014015   0.17707638119406133   0.3959760865280266   0.5503463238379555   0.8847575653255588   0.05281955579777341   0.3531733722649761   0.10696237348267852   0.6351079899268456   0.7880708786742354   0.1367988332000336   0.7386245470747731   0.5240071356561498   0.6490949618163243   0.8332348076034916   0.06039986005936   0.6075311125258632   0.9914556119908984   0.8575098402968061   0.7691887804586959   0.5444757412793814   0.2358361539220206   0.5855343707475156   0.8201351006606037   0.23670692010924127   0.05875977272795925   0.18955828421948898   0.26978877682264824   0.3519493547836825   0.0059402169301858414   0.8363849119545129   0.1628264033399697   0.7168413648568369   0.21786933825595045   0.6995860787544793   0.42420185626519663   0.1928342292006871   0.5687743764396261   0.8663512711509876   0.36380199620583664   0.5853031166748238   0.5773187644487278   0.008841430854181534   0.5946132157471408   0.04082737539544245   0.34148261052670714   0.4233070601066659   0.7744781150865371   0.8041204552862011   0.2827228377987479   0.23374877588717693   0.5046893382638888   0.4521711005025187   0.27678262086856203   0.39736386393266404   0.3418629349239191   0.7353297356456818   0.058913282612611605   0.6977777851781848   0.9176610786587225   0.5424955064449948   0.4901389061729855   0.8314265140271971
0.5538590824528858   0.9571923897701708   0.9128201417242577   0.8225850831730156   0.9592458667057452   0.9163650143747284   0.5713375311975506   0.3992780230663497   0.1847677516192081   0.11224455908852723   0.28861469339880275   0.16552924717917272   0.6800784133553193   0.6600734585860085   0.011832072530240698   0.7681653832465086   0.33821547843140015   0.9247437229403267   0.9529187899176291   0.07038759806832386   0.4205543997726776   0.382248216495332   0.46277988374464357   0.23896108404112673   0.8666953173197918   0.4250558267251611   0.5499597420203858   0.41637600086811116   0.9074494506140466   0.5086908123504328   0.9786222108228352   0.0170979778017615   0.7226816989948385   0.3964462532619055   0.6900075174240324   0.8515687306225888   0.04260328563951922   0.736372794675897   0.6781754448937917   0.08340334737608014   0.7043878072081191   0.8116290717355702   0.7252566549761625   0.013015749307756291   0.2838334074354415   0.4293808552402382   0.262476771231519   0.7740546652666296   0.41713809011564973   0.004325028515077065   0.7125170292111332   0.35767866439851836   0.5096886395016031   0.4956342161646443   0.7338948183882981   0.3405806865967569   0.7870069405067647   0.09918796290273883   0.04388730096426572   0.4890119559741681   0.7444036548672455   0.3628151682268419   0.365711856070474   0.40560860859808795
0.04001584765912638   0.5511860964912717   0.6404552010943114   0.39259285929033166   0.7561824402236849   0.12180524125103347   0.37797842986279245   0.6185381940237021   0.33904435010803513   0.1174802127359564   0.6654614006516592   0.2608595296251837   0.829355710606432   0.621845996571312   0.9315665822633611   0.9202788430284269   0.0423487700996673   0.5226580336685732   0.8876792812990953   0.43126688705425875   0.29794511523242184   0.15984286544173135   0.5219674252286213   0.025658278456170774   0.2579292675732955   0.6086567689504597   0.8815122241343099   0.6330654191658391   0.5017468273496105   0.48685152769942625   0.5035337942715175   0.014527225142136991   0.1627024772415754   0.3693713149634698   0.8380723936198583   0.7536676955169532   0.3333467666351434   0.7475253183921577   0.9065058113564972   0.8333888524885265   0.2909979965354761   0.22486728472358453   0.0188265300574018   0.4021219654342677   0.9930528813030542   0.06502441928185318   0.4968591048287805   0.3764636869780969   0.7351236137297588   0.4563676503313935   0.6153468806944706   0.7433982678122578   0.23337678638014825   0.9695161226319673   0.11181308642295314   0.7288710426701208   0.07067430913857284   0.6001448076684974   0.2737406928030949   0.9752033471531676   0.7373275425034295   0.8526194892763397   0.3672348814465977   0.14181449466464113
0.4463295459679533   0.6277522045527552   0.3484083513891959   0.7396925292303734   0.453276664664899   0.562727785270902   0.8515492465604154   0.36322884225227653   0.7181530509351403   0.10636013493950848   0.23620236586594487   0.6198305744400187   0.484776264554992   0.1368440123075412   0.12438927944299172   0.8909595317698978   0.41410195541641914   0.5366992046390437   0.8506485866398968   0.9157561846167304   0.6767744129129897   0.6840797153627041   0.4834137051932991   0.7739416899520892   0.2304448669450364   0.05632751080994891   0.1350053538041032   0.03424916072171576   0.7771682022801374   0.4935997255390469   0.28345610724368775   0.6710203184694392   0.05901515134499712   0.38723959059953844   0.04725374137774289   0.051189744029420545   0.5742388867900051   0.25039557829199727   0.9228644619347511   0.16023021225952266   0.160136931373586   0.7136963736529535   0.07221587529485433   0.24447402764279236   0.4833625184605963   0.029616658290249422   0.5888021701015552   0.4705323376907032   0.2529176515155599   0.9732891474803005   0.453796816297452   0.4362831769689874   0.4757494492354225   0.4796894219412536   0.17034070905376428   0.7652628584995481   0.41673429789042543   0.09244983134171512   0.12308696767602138   0.7140731144701277   0.8424954111004203   0.8420542530497179   0.2002225057412702   0.553842902210605
0.6823584797268343   0.12835787939676438   0.1280066304464159   0.3093688745678126   0.198995961266238   0.09874122110651497   0.5392044603448607   0.8388365368771095   0.9460783097506781   0.12545207362621447   0.08540764404740865   0.402553359908122   0.4703288605152556   0.6457626516849608   0.9150669349936444   0.6372905014085738   0.053594562624830165   0.5533128203432458   0.791979967317623   0.9232173869384462   0.2110991515244099   0.7112585672935279   0.5917574615763528   0.3693744847278413   0.5287406717975757   0.5829006878967635   0.4637508311299369   0.060005610160028686   0.32974471053133764   0.4841594667902485   0.9245463707850763   0.22116907328291927   0.3836664007806595   0.35870739316403405   0.8391387267376675   0.8186157133747972   0.9133375402654039   0.7129447414790732   0.9240717917440232   0.1813252119662234   0.8597429776405737   0.15963192113582744   0.1320918244264002   0.2581078250277772   0.6486438261161639   0.44837335384229954   0.5403343628500474   0.8887333402999359   0.11990315431858826   0.8654726659455361   0.07658353172011048   0.8287277301399072   0.7901584437872506   0.38131319915528755   0.15203716093503425   0.607558656856988   0.40649204300659114   0.02260580599125346   0.3128984341973667   0.7889429434821907   0.49315450274118716   0.3096610645121803   0.3888266424533435   0.6076177315159673
0.6334115251006134   0.15002914337635284   0.2567348180269433   0.34950990648819014   0.9847676989844495   0.7016557895340533   0.7164004551768959   0.46077656618825424   0.8648645446658613   0.8361831235885172   0.6398169234567854   0.632048836048347   0.07470610087861063   0.45486992443322966   0.4877797625217512   0.024490179191359065   0.6682140578720195   0.4322641184419762   0.17488132832438452   0.23554723570916836   0.1750595551308323   0.12260305392979594   0.7860546858710411   0.627929504193201   0.5416480300302189   0.9725739105534431   0.5293198678440978   0.27841959770501096   0.5568803310457694   0.27091812101938983   0.8129194126672019   0.8176430315167568   0.6920157863799081   0.4347349974308726   0.17310248921041646   0.18559419546840972   0.6173096855012975   0.9798650729976429   0.6853227266886652   0.16110401627705065   0.949095627629278   0.5476009545556667   0.5104413983642807   0.9255567805678823   0.7740360724984456   0.4249979006258708   0.7243867124932397   0.2976272763746812   0.23238804246822678   0.4524239900724277   0.1950668446491419   0.019207678669670256   0.6755077114224575   0.18150586905303787   0.38214743198194   0.20156464715291353   0.9834919250425493   0.7467708716221653   0.20904494277152355   0.015970451684503808   0.36618223954125184   0.7669057986245222   0.5237222160828583   0.8548664354074531
0.4170866119119739   0.21930484406885553   0.013280817718577568   0.9293096548395708   0.6430505394135282   0.7943069434429847   0.28889410522533787   0.6316823784648896   0.41066249694530144   0.341882953370557   0.093827260576196   0.6124746997952194   0.735154785522844   0.16037708431751918   0.711679828594256   0.4109100526423059   0.7516628604802946   0.41360621269535397   0.5026348858227324   0.39493960095780206   0.38548062093904284   0.6467004140708317   0.9789126697398741   0.5400731655503489   0.968394009027069   0.42739557000197614   0.9656318520212965   0.6107635107107781   0.32534346961354077   0.6330886265589915   0.6767377467959587   0.9790811322458883   0.9146809726682393   0.2912056731884344   0.5829104862197626   0.366606432450669   0.17952618714539537   0.13082858887091522   0.8712306576255067   0.9556963798083631   0.4278633266651007   0.7172223761755613   0.36859577180277425   0.560756778850561   0.042382705726057866   0.07052196210472961   0.38968310206290013   0.02068361330021209   0.0739886966989889   0.6431263921027535   0.42405125004160354   0.40992010258943407   0.7486452270854481   0.010037765543762036   0.7473135032456449   0.4308389703435457   0.8339642544172088   0.7188320923553276   0.16440301702588223   0.06423253789287671   0.6544380672718134   0.5880035034844124   0.29317235940037556   0.10853615808451363
0.22657474060671268   0.8707811273088512   0.9245765875976013   0.5477793792339526   0.18419203488065483   0.8002591652041215   0.5348934855347012   0.5270957659337405   0.11020333818166592   0.15713277310136808   0.11084223549309768   0.11717566334430647   0.36155811109621777   0.14709500755760604   0.3635287322474528   0.6863366930007608   0.527593856679009   0.4282629152022784   0.19912571522157058   0.6221041551078841   0.8731557894071956   0.840259411717866   0.905953355821195   0.5135679970233705   0.646581048800483   0.9694782844090148   0.9813767682235937   0.9657886177894178   0.4623890139198281   0.1692191192048933   0.4464832826888924   0.43869285185567736   0.35218567573816223   0.012086346103525207   0.33564104719579474   0.32151718851137084   0.9906275646419445   0.8649913385459191   0.9721123149483419   0.6351804955106101   0.4630337079629354   0.43672842334364076   0.7729865997267714   0.01307634040272596   0.5898779185557398   0.5964690116257748   0.8670332439055763   0.49950834337935546   0.9432968697552567   0.62699072721676   0.8856564756819827   0.5337197255899376   0.48090785583542867   0.45777160801186667   0.43917319299309027   0.09502687373426028   0.1287221800972664   0.44568526190834146   0.10353214579729553   0.7735096852228894   0.13809461545532198   0.5806939233624223   0.1314198308489536   0.13832918971227934
0.6750609074923866   0.14396550001878153   0.35843323112218217   0.12525284930955338   0.08518298893664686   0.5474964883930068   0.4913999872166058   0.6257445059301979   0.14188611918139007   0.9205057611762468   0.6057435115346231   0.09202478034026028   0.6609782633459614   0.46273415316438016   0.1665703185415328   0.996997906606   0.532256083248695   0.017048891256038732   0.06303817274423729   0.2234882213831106   0.394161467793373   0.43635496789361644   0.9316183418952837   0.08515903167083128   0.7191005603009865   0.29238946787483494   0.5731851107731015   0.9599061823612779   0.6339175713643396   0.7448929794818282   0.0817851235564957   0.33416167643108   0.49203145218294947   0.8243872183055814   0.4760416120218726   0.24213689609081973   0.8310531888369881   0.3616530651412012   0.3094712934803398   0.2451389894848197   0.29879710558829303   0.34460417388516246   0.2464331207361025   0.021650768101709093   0.9046356377949201   0.908249205991546   0.3148147788408188   0.9364917364308778   0.18553507749393358   0.615859738116711   0.7416296680677174   0.9765855540695999   0.551617506129594   0.8709667586348829   0.6598445445112217   0.6424238776385199   0.05958605394664453   0.04657954032930153   0.183802932489349   0.4002869815477002   0.22853286510965648   0.6849264751881003   0.8743316390090092   0.1551479920628805
0.9297357595213634   0.3403223013029379   0.6278985182729068   0.1334972239611714   0.02510012172644342   0.4320730953113919   0.3130837394320879   0.19700548753029357   0.8395650442325099   0.8162133571946808   0.5714540713643707   0.22041993346069366   0.2879475381029158   0.945246598559798   0.911609526853149   0.5779960558221737   0.22836148415627128   0.8986670582304964   0.7278065943638   0.17770907427447352   0.9998286190466148   0.21374058304239604   0.8534749553547908   0.022561082211593038   0.07009285952525139   0.8734182817394581   0.22557643708188407   0.8890638582504217   0.04499273779880797   0.44134518642806625   0.9124926976497961   0.6920583707201281   0.20542769356629814   0.6251318292333854   0.34103862628542553   0.4716384372594344   0.9174801554633824   0.6798852306735875   0.42942909943227653   0.8936423814372607   0.689118671307111   0.7812181724430911   0.7016225050684765   0.7159333071627871   0.6892900522604962   0.567477589400695   0.8481475497136857   0.6933722249511941   0.6191971927352449   0.6940593076612369   0.6225711126318016   0.8043083667007724   0.5742044549364369   0.25271412123317066   0.7100784149820055   0.1122499959806444   0.3687767613701387   0.6275822919997852   0.36903978869658   0.64061155872121   0.4512966059067564   0.9476970613261977   0.9396106892643035   0.7469691772839493
0.7621779345996453   0.16647888888310663   0.23798818419582699   0.031035870121162185   0.07288788233914915   0.5990012994824115   0.3898406344821413   0.3376636451699681   0.45369068960390435   0.9049419918211746   0.7672695218503396   0.5333552784691956   0.8794862346674674   0.6522278705880039   0.05719110686833413   0.4211052824885512   0.5107094732973287   0.02464557858821872   0.6881513181717541   0.7804937237673412   0.05941286739057234   0.07694851726202098   0.7485406289074507   0.03352454648339189   0.29723493279092694   0.9104696283789143   0.5105524447116236   0.0024886763622297076   0.2243470504517778   0.31146832889650283   0.12071181022948241   0.6648250311922617   0.7706563608478735   0.4065263370753282   0.35344228837914277   0.13146975272306602   0.891170126180406   0.7542984664873242   0.29625118151080865   0.7103644702345148   0.3804606528830773   0.7296528878991055   0.6080998633390545   0.9298707464671736   0.32104778549250496   0.6527043706370845   0.8595592344316039   0.8963461999837817   0.02381285270157797   0.7422347422581701   0.3490067897199801   0.893857523621552   0.7994658022498001   0.4307664133616673   0.22829497949049773   0.22903249242929036   0.02880944140192668   0.02424007628633917   0.874852691111355   0.09756273970622435   0.13763931522152067   0.26994160979901494   0.5786015096005463   0.38719826947170954
0.7571786623384434   0.5402887218999095   0.9705016462614918   0.45732752300453594   0.4361308768459385   0.887584351262825   0.11094241182988798   0.5609813230207543   0.4123180241443605   0.1453496090046548   0.7619356221099078   0.6671237993992023   0.6128522218945603   0.7145831956429874   0.5336406426194101   0.43809130696991194   0.5840427804926337   0.6903431193566483   0.6587879515080551   0.3405285672636876   0.44640346527111296   0.42040150955763333   0.08018644190750887   0.953330297791978   0.6892248029326696   0.8801127876577238   0.10968479564601707   0.4960027747874421   0.25309392608673115   0.992528436394899   0.9987423838161291   0.9350214517666878   0.8407759019423706   0.8471788273902441   0.23680676170622122   0.26789765236748553   0.2279236800478103   0.1325956317472567   0.7031661190868111   0.8298063453975736   0.6438808995551767   0.4422525123906084   0.044378167578755935   0.489277778133886   0.19747743428406367   0.021851002832975086   0.9641917256712471   0.535947480341908   0.5082526313513941   0.14173821517525123   0.85450693002523   0.03994470555446593   0.25515870526466294   0.1492097787803523   0.8557645462091009   0.10492325378777813   0.4143828033222923   0.30203095139010816   0.6189577845028796   0.8370256014202926   0.186459123274482   0.1694353196428515   0.9157916654160686   0.00721925602271901
0.5425782237193053   0.727182807252243   0.8714134978373126   0.5179414778888329   0.3451007894352417   0.705331804419268   0.9072217721660656   0.981993997546925   0.8368481580838476   0.5635935892440168   0.052714842140835556   0.942049291992459   0.5816894528191847   0.41438381046366446   0.19695029593173466   0.8371260382046809   0.1673066494968924   0.1123528590735563   0.577992511428855   0.00010043678438833529   0.9808475262224103   0.9429175394307048   0.6622008460127864   0.9928811807616693   0.43826930250310503   0.2157347321784617   0.7907873481754738   0.4749397028728363   0.09316851306786332   0.5104029277591937   0.8835655760094082   0.49294570532591137   0.2563203549840157   0.9468093385151769   0.8308507338685727   0.5508964133334523   0.674630902164831   0.5324255280515124   0.633900437936838   0.7137703751287713   0.5073242526679386   0.42007266897795614   0.05590792650798307   0.713669938344383   0.5264767264455282   0.47715512954725137   0.39370708049519665   0.7207887575827137   0.08820742394242317   0.26142039736878964   0.6029197323197228   0.24584905470987733   0.9950389108745599   0.7510174696095959   0.7193541563103145   0.752903349383966   0.7387185558905441   0.804208131094419   0.8885034224417419   0.20200693605051373   0.0640876537257132   0.2717826030429066   0.25460298450490376   0.4882365609217424
0.5567634010577747   0.8517099340649504   0.1986950579969207   0.7745666225773594   0.030286674612246423   0.37455480451769907   0.804987977501724   0.05377786499464572   0.9420792506698232   0.11313440714890943   0.20206824518200125   0.8079288102847684   0.9470403397952634   0.3621169375393135   0.4827140888716867   0.055025460900802396   0.2083217839047192   0.5579088064448945   0.5942106664299449   0.8530185248502887   0.144234130179006   0.28612620340198797   0.3396076819250411   0.3647819639285463   0.5874707291212313   0.43441626933703753   0.14091262392812043   0.5902153413511869   0.5571840545089849   0.05986146481933848   0.33592464642639636   0.5364374763565412   0.6151048038391617   0.9467270576704291   0.13385640124439507   0.7285086660717728   0.6680644640438983   0.5846101201311156   0.6511423123727084   0.6734832051709704   0.4597426801391791   0.026701313686221032   0.05693164594276348   0.8204646803206818   0.31550854996017313   0.7405751102842331   0.7173239640177224   0.4556827163921354   0.7280378208389418   0.30615884094719553   0.5764113400896019   0.8654673750409485   0.17085376632995686   0.24629737612785707   0.2404866936632056   0.32902989868440735   0.5557489624907952   0.299570318457428   0.1066302924188105   0.6005212326126346   0.8876844984468969   0.7149601983263125   0.45548798004610214   0.9270380274416642
0.42794181830771777   0.6882588846400914   0.3985563341033387   0.10657334712098245   0.11243326834754462   0.9476837743558584   0.6812323700856163   0.650890630728847   0.3843954475086028   0.6415249334086628   0.10482102999601436   0.7854232556878985   0.213541681178646   0.3952275572808058   0.8643343363328088   0.4563933570034912   0.6577927186878508   0.09565723882337775   0.7577040439139983   0.8558721243908567   0.7701082202409539   0.38069704049706526   0.3022160638678961   0.9288340969491925   0.3421664019332362   0.6924381558569739   0.9036597297645574   0.8222607498282101   0.22973313358569158   0.7447543815011155   0.22242735967894114   0.17137011909936303   0.8453376860770887   0.10322944809245266   0.1176063296829268   0.3859468634114645   0.6317960048984428   0.7080018908116469   0.253271993350118   0.9295535064079733   0.974003286210592   0.6123446519882692   0.49556794943611976   0.07368138201711669   0.203895065969638   0.2316476114912039   0.19335188556822366   0.1448472850679242   0.8617286640364018   0.5392094556342301   0.2896921558036662   0.32258653523971415   0.6319955304507102   0.7944550741331146   0.06726479612472505   0.15121641614035114   0.7866578443736214   0.691225626040662   0.9496584664417983   0.7652695527288866   0.15486183947517868   0.983223735229015   0.6963864730916802   0.8357160463209133
0.18085855326458672   0.37087908324074587   0.20081852365556047   0.7620346643037966   0.9769634872949488   0.13923147174954198   0.007466638087336814   0.6171873792358724   0.11523482325854692   0.6000220161153119   0.7177744822836706   0.29460084399615827   0.48323929280783673   0.8055669419821974   0.6505096861589456   0.14338442785580713   0.6965814484342153   0.11434131594153546   0.7008512197171473   0.3781148751269205   0.5417196089590366   0.13111758071252044   0.004464746625467063   0.5423988288060072   0.36086105569444993   0.7602384974717746   0.8036462229699066   0.7803641645022106   0.3838975683995012   0.6210070257222327   0.7961795848825698   0.16317678526633816   0.2686627451409543   0.020985009606920697   0.07840510259889917   0.8685759412701799   0.7854234523331175   0.21541806762472335   0.4278954164399536   0.7251915134143727   0.08884200389890225   0.10107675168318789   0.7270441967228063   0.3470766382874523   0.5471223949398656   0.9699591709706674   0.7225794500973393   0.8046778094814451   0.1862613392454157   0.20972067349889284   0.9189332271274326   0.02431364497923445   0.8023637708459145   0.5887136477766602   0.12275364224486286   0.8611368597128963   0.5337010257049603   0.5677286381697395   0.0443485396459637   0.9925609184427163   0.7482775733718428   0.3523105705450162   0.6164531232060101   0.2673694050283436
0.6594355694729405   0.25123381886182833   0.8894089264832038   0.9202927667408913   0.11231317453307488   0.28127464789116086   0.16682947638586454   0.11561495725944632   0.9260518352876591   0.07155397439226803   0.2478962492584319   0.09130131228021186   0.12368806444174463   0.48284032661560783   0.12514260701356905   0.2301644525673156   0.5899870387367844   0.9151116884458683   0.08079406736760535   0.23760353412459922   0.8417094653649416   0.5628011179008521   0.46434094416159527   0.9702341290962556   0.18227389589200113   0.3115672990390238   0.5749320176783914   0.049941362355364234   0.06996072135892625   0.030292651147862944   0.4081025412925269   0.9343264050959179   0.1439088860712671   0.9587386767555949   0.160206292034095   0.843025092815706   0.020220821629522465   0.4758983501399871   0.03506368502052596   0.6128606402483905   0.4302337828927381   0.5607866616941188   0.9542696176529206   0.37525710612379126   0.5885243175277964   0.9979855437932666   0.48992867349132535   0.40502297702753565   0.4062504216357954   0.6864182447542428   0.9149966558129339   0.3550816146721714   0.3362897002768691   0.6561255936063799   0.506894114520407   0.4207552095762535   0.19238081420560205   0.697386916850785   0.346687822486312   0.5777301167605474   0.17215999257607956   0.22148856671079792   0.31162413746578604   0.9648694765121569
0.7419262096833414   0.6607019050166791   0.3573545198128654   0.5896123703883658   0.15340189215554498   0.6627163612234124   0.8674258463215401   0.18458939336083008   0.7471514705197496   0.9762981164691695   0.9524291905086062   0.8295077786886587   0.41086177024288045   0.32017252286278963   0.44553507598819914   0.40875256911240515   0.21848095603727843   0.6227856060120046   0.09884725350188713   0.8310224523518577   0.04632096346119887   0.4012970393012067   0.7872231160361011   0.8661529758397007   0.3043947537778574   0.7405951342845276   0.42986859622323564   0.276540605451335   0.15099286162231243   0.07787877306111514   0.5624427499016955   0.09195121209050493   0.40384139110256284   0.1015806565919456   0.6100135593930894   0.2624434334018463   0.9929796208596824   0.781408133729156   0.16447848340489027   0.8536908642894411   0.7744986648224039   0.15862252771715135   0.06563122990300316   0.022668411937583365   0.7281777013612051   0.7573254884159446   0.2784081138669021   0.15651543609788263   0.42378294758334767   0.016730354131417078   0.8485395176436664   0.8799748306465476   0.2727900859610352   0.938851581070302   0.2860967677419709   0.7880236185560426   0.8689486948584724   0.8372709244783564   0.6760832083488815   0.5255801851541965   0.87596907399879   0.055862790749200385   0.5116047249439912   0.6718893208647553
0.10147040917638608   0.8972402630320491   0.44597349504098804   0.649220908927172   0.37329270781518104   0.13991477461610438   0.16756538117408598   0.49270547282928934   0.9495097602318334   0.1231844204846873   0.3190258635304195   0.6127306421827418   0.6767196742707982   0.18433283941438536   0.0329290957884486   0.824707023626699   0.8077709794123258   0.347061914936029   0.35684588743956713   0.29912683847250265   0.9318019054135358   0.29119912418682864   0.8452411624955759   0.6272375176077473   0.8303314962371497   0.3939588611547796   0.3992676674545878   0.9780166086805754   0.45703878842196866   0.2540440865386752   0.23170228628050185   0.485311135851286   0.5075290281901353   0.13085966605398794   0.9126764227500823   0.8725804936685443   0.8308093539193371   0.9465268266396025   0.8797473269616337   0.04787347004184521   0.02303837450701134   0.5994649117035735   0.5229014395220667   0.7487466315693425   0.09123646909347556   0.3082657875167449   0.6776602770264908   0.12150911396159526   0.26090497285632586   0.9143069263619653   0.2783926095719029   0.14349250528101992   0.8038661844343572   0.66026283982329   0.046690323291401076   0.6581813694297339   0.2963371562442219   0.5294031737693021   0.1340139005413187   0.7856008757611896   0.4655278023248848   0.5828763471296996   0.25426657357968496   0.7377274057193445
0.4424894278178734   0.9834114354261261   0.7313651340576183   0.9889807741500019   0.3512529587243979   0.6751456479093811   0.05370485703112752   0.8674716601884066   0.09034798586807201   0.7608387215474158   0.7753122474592246   0.7239791549073867   0.2864818014337148   0.10057588172412575   0.7286219241678236   0.06579778547765279   0.990144645189493   0.5711727079548236   0.5946080236265048   0.28019690971646316   0.5246168428646082   0.9882963608251241   0.34034145004681987   0.5424695039971187   0.08212741504673475   0.004884925398997973   0.6089763159892015   0.5534887298471168   0.7308744563223369   0.32973927748961684   0.5552714589580741   0.6860170696587102   0.6405264704542649   0.568900555942201   0.7799592114988495   0.9620379147513235   0.35404466902055004   0.4683246742180753   0.05133728733102595   0.8962401292736707   0.36390002383105713   0.8971519662632517   0.45672926370452116   0.6160432195572075   0.8392831809664489   0.9088556054381276   0.11638781365770129   0.07357371556008888   0.7571557659197142   0.9039706800391296   0.5074114976684997   0.520084985712972   0.026281309597377314   0.5742314025495129   0.9521400387104256   0.8340679160542619   0.3857548391431124   0.005330846607311821   0.1721808272115762   0.8720300013029384   0.031710170122562366   0.5370061723892365   0.12084353988055027   0.9757898720292677
0.6678101462915053   0.6398542061259849   0.6641142761760291   0.35974665247206006   0.8285269653250563   0.7309986006878573   0.5477264625183278   0.2861729369119712   0.07137119940534209   0.8270279206487277   0.0403149648498281   0.7660879511989991   0.04508988980796477   0.2527965180992148   0.08817492613940241   0.9320200351447373   0.6593350506648523   0.24746567149190296   0.9159940989278262   0.05999003384179891   0.6276248805422899   0.7104594991026664   0.7951505590472759   0.08420016181253126   0.9598147342507848   0.07060529297668149   0.1310362828712468   0.7244535093404711   0.13128776892572844   0.33960669228882423   0.583309820352919   0.4382805724285   0.05991656952038636   0.5125787716400966   0.5429948555030909   0.6721926212295009   0.014826679712421591   0.2597822535408818   0.4548199293636885   0.7401725860847636   0.35549162904756926   0.012316582048978857   0.5388258304358623   0.6801825522429646   0.7278667485052793   0.30185708294631247   0.7436752713885864   0.5959823904304334   0.7680520142544945   0.23125178996963097   0.6126389885173396   0.8715288810899622   0.6367642453287661   0.8916450976808068   0.029329168164420574   0.43324830866146224   0.5768476758083797   0.37906632604071017   0.4863343126613297   0.7610556874319614   0.5620209960959581   0.11928407249982836   0.03151438329764123   0.020883101347197765
0.2065293670483889   0.10696749045084951   0.492688552861779   0.3407005491042331   0.4786626185431096   0.805110407504537   0.7490132814731926   0.7447181586737996   0.7106106042886151   0.5738586175349061   0.13637429295585307   0.8731892775838375   0.07384635895984898   0.6822135198540993   0.10704512479143248   0.4399409689223752   0.4969986831514692   0.3031471938133891   0.6207108121301028   0.6788852814904138   0.9349776870555111   0.18386312131356072   0.5891964288324616   0.6580021801432161   0.7284483200071222   0.07689563086271123   0.0965078759706826   0.317301631038983   0.2497857014640126   0.2717852233581742   0.34749459449749   0.5725834723651834   0.5391750971753975   0.6979266058232682   0.2111203015416369   0.6993941947813459   0.46532873821554854   0.01571308596916885   0.10407517675020445   0.25945322585897074   0.9683300550640793   0.7125658921557797   0.4833643646201016   0.5805679443685569   0.03335236800856819   0.5287027708422191   0.8941679357876401   0.9225657642253409   0.304904048001446   0.4518071399795078   0.7976600598169575   0.6052641331863579   0.05511834653743338   0.1800219166213336   0.4501654653194675   0.032680660821174504   0.5159432493620358   0.48209531079806545   0.23904516377783058   0.3332864660398286   0.05061451114648732   0.46638222482889663   0.13496998702762614   0.07383324018085789
0.08228445608240803   0.7538163326731169   0.6516056224075245   0.493265295812301   0.04893208807383984   0.22511356183089784   0.7574376866198844   0.5706995315869602   0.7440280400723939   0.7733064218513901   0.9597776268029269   0.9654353984006023   0.6889096935349605   0.5932845052300565   0.5096121614834593   0.9327547375794278   0.17296644417292462   0.111189194431991   0.2705669977056288   0.5994682715395993   0.12235193302643729   0.6448069696030944   0.13559701067800264   0.5256350313587413   0.04006747694402926   0.8909906369299775   0.48399138827047816   0.03236973554644036   0.9911353888701894   0.6658770750990797   0.7265537016505937   0.46167020395948016   0.24710734879779556   0.8925706532476896   0.7667760748476669   0.49623480555887783   0.558197655262835   0.29928614801763315   0.25716391336420746   0.5634800679794499   0.38523121108991043   0.18809695358564213   0.9865969156585787   0.9640117964398507   0.26287927806347317   0.5432899839825478   0.8509999049805761   0.43837676508110934   0.2228118011194439   0.6522993470525702   0.36700851671009793   0.406007029534669   0.23167641224925448   0.9864222719534905   0.6404548150595042   0.9443368255751888   0.9845690634514589   0.0938516187058009   0.8736787402118373   0.448102020016311   0.42637140818862385   0.7945654706881677   0.6165148268476298   0.884621952036861
0.0411401970987134   0.6064685171025256   0.6299179111890512   0.9206101555970103   0.7782609190352402   0.06317853311997786   0.7789180062084752   0.4822333905159009   0.5554491179157963   0.41087918606740764   0.41190948949837725   0.07622636098123195   0.32377270566654187   0.4244569141139171   0.7714546744388731   0.13188953540604312   0.339203642215083   0.33060529540811623   0.8977759342270357   0.6837875153897321   0.9128322340264591   0.5360398247199485   0.28126110737940585   0.7991655633528711   0.8716920369277457   0.9295713076174229   0.6513431961903546   0.8785554077558608   0.09343111789250544   0.866392774497445   0.8724251899818796   0.39632201723995986   0.537981999976709   0.45551358843003736   0.4605157004835023   0.32009565625872793   0.21420929431016722   0.03105667431612025   0.6890610260446293   0.1882061208526848   0.8750056520950843   0.700451378908004   0.7912850918175935   0.5044186054629527   0.9621734180686251   0.16441155418805553   0.5100239844381876   0.7052530421100816   0.09048138114087946   0.23484024657063265   0.858680788247833   0.8266976343542207   0.997050263248374   0.3684474720731876   0.9862555982659534   0.4303756171142609   0.45906826327166494   0.9129338836431502   0.5257398977824511   0.11027996085553299   0.24485896896149772   0.88187720932703   0.8366788717378218   0.9220738400028482
0.3698533168664135   0.18142583041902596   0.04539377992022836   0.41765523453989556   0.4076798987977883   0.01701427623097044   0.5353697954820407   0.712402192429814   0.3171985176569089   0.7821740296603378   0.6766890072342077   0.8857045580755932   0.32014825440853484   0.41372655758715016   0.6904334089682542   0.4553289409613323   0.86107999113687   0.500792673944   0.1646935111858031   0.3450489801057993   0.6162210221753722   0.6189154646169699   0.3280146394479812   0.4229751401029511   0.24636770530895874   0.43748963419794396   0.28262085952775284   0.005319905563055587   0.8386878065111705   0.42047535796697355   0.7472510640457122   0.2929177131332416   0.5214892888542616   0.6383013283066358   0.07056205681150444   0.40721315505764843   0.20134103444572676   0.22457477071948556   0.3801286478432502   0.9518842140963161   0.3402610433088568   0.7237820967754857   0.2154351366574471   0.6068352339905168   0.7240400211334846   0.1048666321585157   0.8874204972094659   0.18386009388756566   0.4776723158245259   0.6673769979605717   0.604799637681713   0.17854018832451007   0.6389845093133555   0.2469016399935982   0.8575485736360009   0.8856224751912685   0.11749522045909386   0.6086003116869625   0.7869865168244964   0.47840932013362003   0.9161541860133671   0.3840255409674769   0.4068578689812462   0.526525106037304
0.5758931427045103   0.6602434441919912   0.1914227323237991   0.9196898720467872   0.8518531215710257   0.5553768120334756   0.3040022351143333   0.7358297781592215   0.37418080574649976   0.8879998140729038   0.6992025974326203   0.5572895898347114   0.7351962964331443   0.6410981740793056   0.8416540237966194   0.671667114643443   0.6177010759740504   0.03249786239234314   0.05466750697212298   0.1932577945098229   0.7015468899606834   0.6484723214248662   0.6478096379908768   0.666732688472519   0.12565374725617307   0.988228877232875   0.4563869056670777   0.7470428164257318   0.27380062568514746   0.43285206519939945   0.1523846705527444   0.011213038266510298   0.8996198199386477   0.5448522511264957   0.45318207312012415   0.4539234484317989   0.16442352350550343   0.90375407704719   0.6115280493235048   0.7822563337883559   0.546722447531453   0.8712562146548469   0.5568605423513818   0.5889985392785331   0.8451755575707697   0.22278389322998068   0.9090509043605051   0.9222658508060141   0.7195218103145966   0.23455501599710565   0.4526639986934274   0.1752230343802823   0.44572118462944915   0.8017029507977061   0.300279328140683   0.164009996113772   0.5461013646908014   0.25685069967121055   0.8470972550205588   0.7100865476819731   0.38167784118529796   0.3530966226240205   0.23556920569705403   0.9278302138936172
0.834955393653845   0.48184040796917355   0.6787086633456723   0.3388316746150841   0.9897798360830753   0.2590565147391929   0.7696577589851672   0.41656582380907003   0.27025802576847874   0.02450149874208721   0.31699376029173976   0.24134278942878773   0.8245368411390296   0.222798547944381   0.0167144321510568   0.07733279331501572   0.2784354764482282   0.9659478482731705   0.16961717713049798   0.3672462456330426   0.8967576352629302   0.61285122564915   0.934047971433444   0.43941603173942545   0.06180224160908523   0.13101081767997644   0.2553393080877718   0.10058435712434129   0.07202240552600991   0.8719543029407836   0.4856815491026046   0.6840185333152713   0.8017643797575312   0.8474528041986964   0.1686877888108648   0.4426757438864835   0.9772275386185016   0.6246542562543154   0.151973356659808   0.3653429505714678   0.6987920621702735   0.6587064079811449   0.98235617952931   0.9980967049384252   0.8020344269073433   0.04585518233199488   0.04830820809586605   0.5586806731989997   0.740232185298258   0.9148443646520185   0.7929689000080943   0.4580963160746585   0.668209779772248   0.042890061711234856   0.3072873509054897   0.7740777827593872   0.8664454000147169   0.1954372575125385   0.13859956209462493   0.3314020388729037   0.8892178613962153   0.5707830012582231   0.9866262054348169   0.9660590883014359
0.19042579922594183   0.9120765932770782   0.004270025905506909   0.9679623833630108   0.3883913723185986   0.8662214109450834   0.9559618178096408   0.40928171016401094   0.6481591870203406   0.951377046293065   0.16299291780154657   0.9511853940893524   0.9799494072480925   0.9084869845818301   0.8557055668960568   0.17710761132996525   0.11350400723337559   0.7130497270692916   0.7171060048014319   0.8457055724570616   0.2242861458371603   0.14226672581106847   0.730479799366615   0.8796464841556256   0.03386034661121848   0.2301901325339902   0.726209773461108   0.9116841007926149   0.6454689742926198   0.3639687215889068   0.7702479556514672   0.5024023906286039   0.9973097872722793   0.41259167529584184   0.6072550378499206   0.5512169965392515   0.01736038002418681   0.5041046907140118   0.7515494709538638   0.3741093852092862   0.9038563727908112   0.7910549636447202   0.034443466152431906   0.5284038127522247   0.6795702269536509   0.6487882378336517   0.30396366678581693   0.6487573285965991   0.6457098803424324   0.41859810529966146   0.5777538933247088   0.7370732278039842   0.0002409060498125479   0.05462938371075466   0.8075059376732416   0.2346708371753802   0.00293111877753325   0.6420377084149128   0.20025089982332092   0.6834538406361288   0.9855707387533464   0.13793301770090108   0.4487014288694571   0.3093444554268425
0.08171436596253522   0.34687805405618094   0.4142579627170252   0.7809406426746178   0.4021441390088843   0.6980898162225293   0.11029429593120828   0.13218331407801878   0.7564342586664519   0.27949171092286784   0.5325404026064995   0.3951100862740346   0.7561933526166393   0.22486232721211316   0.7250344649332578   0.16043924909865442   0.7532622338391061   0.5828246187972004   0.524783565109937   0.4769854084625257   0.7676914950857596   0.44489160109629927   0.07608213624047984   0.16764095303568313   0.6859771291232244   0.09801354704011832   0.6618241735234547   0.3867003103610653   0.2838329901143401   0.39992373081758903   0.5515298775922464   0.2545169962830465   0.5273987314478882   0.1204320198947212   0.01898947498574691   0.8594069100090119   0.7712053788312488   0.895569692682608   0.29395501005248903   0.6989676609103574   0.0179431449921428   0.3127450738854077   0.7691714449425521   0.22198225244783182   0.25025164990638316   0.8678534727891084   0.6930893087020723   0.054341299412148665   0.5642745207831588   0.7698399257489901   0.03126513517861765   0.6676409890510834   0.2804415306688186   0.36991619493140104   0.47973525758637126   0.41312399276803685   0.7530427992209304   0.24948417503667983   0.4607457826006244   0.553717082759025   0.9818374203896815   0.3539144823540718   0.16679077254813532   0.8547494218486675
0.9638942753975387   0.04116940846866413   0.3976193276055832   0.6327671694008357   0.7136426254911555   0.17331593567955572   0.7045300189035109   0.5784258699886871   0.14936810470799683   0.40347600993056565   0.6732648837248932   0.9107848809376037   0.8689265740391782   0.03355981499916461   0.19352962613852198   0.49766088816956683   0.11588377481824784   0.7840756399624847   0.7327838435378976   0.9439438054105418   0.13404635442856636   0.43016115760841295   0.5659930709897623   0.0891943835618743   0.17015207903102766   0.3889917491397488   0.1683737433841791   0.4564272141610386   0.45650945353987216   0.2156758134601931   0.4638437244806682   0.8780013441723515   0.3071413488318753   0.8121998035296274   0.7905788407557749   0.9672164632347479   0.4382147747926971   0.7786399885304628   0.5970492146172529   0.46955557506518103   0.32233099997444925   0.994564348567978   0.8642653710793553   0.5256117696546393   0.18828464554588292   0.5644031909595651   0.29827230008959305   0.4364173860927649   0.01813256651485524   0.17541144181981627   0.12989855670541395   0.9799901719317263   0.5616231129749831   0.9597356283596231   0.6660548322247457   0.10198882775937483   0.2544817641431078   0.14753582482999572   0.8754759914689708   0.134772364524627   0.8162669893504106   0.3688958362995329   0.2784267768517179   0.665216789459446
0.49393598937596145   0.37433148773155484   0.41416140577236255   0.1396050198048067   0.3056513438300785   0.8099282967719897   0.1158891056827695   0.7031876337120417   0.2875187773152233   0.6345168549521735   0.9859905489773556   0.7231974617803154   0.7258956643402401   0.6747812265925504   0.3199357167526098   0.6212086340209405   0.47141390019713236   0.5272454017625546   0.444459725283639   0.4864362694963136   0.6551469108467217   0.1583495654630217   0.16603294843192107   0.8212194800368676   0.16121092147076024   0.7840180777314669   0.7518715426595586   0.681614460232061   0.8555595776406817   0.9740897809594772   0.635982436976789   0.9784268265200192   0.5680408003254585   0.33957292600730365   0.6499918879994335   0.25522936473970387   0.8421451359852183   0.6647916994147534   0.3300561712468237   0.6340207307187633   0.3707312357880859   0.13754629765219875   0.8855964459631848   0.14758446122244975   0.7155843249413643   0.979196732189177   0.7195634975312637   0.3263649811855821   0.554373403470604   0.19517865445771018   0.9676919548717051   0.6447505209535211   0.6988138258299222   0.22108887349823306   0.3317095178949161   0.6663236944335019   0.1307730255044638   0.8815159474909294   0.6817176298954826   0.41109432969379806   0.2886278895192455   0.21672424807617607   0.3516614586486589   0.7770735989750347
0.9178966537311596   0.07917795042397732   0.4660650126854742   0.629489137752585   0.2023123287897953   0.09998121823480027   0.7465015151542106   0.30312415656700287   0.6479389253191913   0.9048025637770901   0.7788095602825055   0.6583736356134817   0.949125099489269   0.6837136902788571   0.4471000423875894   0.9920499411799798   0.8183520739848053   0.8021977427879277   0.7653824124921067   0.5809556114861818   0.5297241844655598   0.5854734947117516   0.41372095384344787   0.8038820125111471   0.6118275307344002   0.5062955442877742   0.9476559411579737   0.1743928747585621   0.40951520194460495   0.406314326052974   0.20115442600376313   0.8712687181915593   0.7615762766254136   0.5015117622758839   0.4223448657212577   0.21289508257807746   0.8124511771361446   0.8177980719970268   0.9752448233336684   0.22084514139809763   0.9940991031513393   0.01560032920909917   0.20986241084156157   0.6398895299119158   0.46437491868577946   0.43012683449734757   0.7961414569981137   0.8360075174007687   0.8525473879513792   0.9238312902095733   0.8484855158401401   0.6616146426422066   0.44303218600677424   0.5175169641565993   0.647331089836377   0.7903459244506474   0.6814559093813606   0.016005201880715404   0.2249862241151193   0.5774508418725699   0.8690047322452161   0.19820712988368858   0.24974140078145096   0.3566057004744723
0.8749056290938768   0.1826068006745894   0.039878989939889385   0.7167161705625565   0.41053071040809735   0.7524799661772418   0.24373753294177566   0.8807086531617878   0.5579833224567181   0.8286486759676686   0.3952520171016356   0.2190940105195811   0.11495113644994387   0.31113171181106924   0.7479209272652586   0.4287480860689337   0.43349522706858323   0.29512650993035383   0.5229347031501393   0.8512972441963638   0.5644904948233671   0.09691938004666527   0.2731933023686884   0.49469154372189145   0.6895848657294903   0.9143125793720759   0.23331431242879902   0.777975373159335   0.279054155321393   0.16183261319483402   0.9895767794870234   0.8972667199975471   0.7210708328646749   0.3331839372271655   0.5943247623853878   0.678172709477966   0.6061196964147311   0.02205222541609625   0.8464038351201292   0.24942462340903235   0.17262446934614778   0.7269257154857424   0.3234691319699898   0.3981273792126686   0.6081339745227806   0.6300063354390771   0.050275829601301385   0.9034358354907772   0.9185491087932903   0.7156937560670013   0.8169615171725023   0.12546046233144226   0.6394949534718973   0.5538611428721673   0.827384737685479   0.2281937423338951   0.9184241206072224   0.22067720564500176   0.23305997530009123   0.5500210328559291   0.3123044241924914   0.1986249802289055   0.3866561401799621   0.3005964094468967
0.1396799548463436   0.4716992647431631   0.06318700820997229   0.9024690302342281   0.5315459803235629   0.8416929293040859   0.012911178608670908   0.999033194743451   0.6129968715302727   0.12599917323708465   0.19594966143616854   0.8735727324120086   0.9735019180583754   0.5721380303649174   0.36856492375068955   0.6453789900781135   0.055077797451152974   0.35146082471991563   0.13550494845059832   0.09535795722218449   0.7427733732586616   0.15283584449101012   0.7488488082706363   0.7947615477752877   0.603093418412318   0.681136579747847   0.685661800060664   0.8922925175410596   0.071547438088755   0.839443650443761   0.672750621451993   0.8932593227976087   0.4585505665584823   0.7134444772066764   0.4768009600158245   0.01968659038560006   0.4850486485001069   0.141306446841759   0.10823603626513496   0.3743076003074865   0.42997085104895394   0.7898456221218434   0.9727310878145367   0.278949643085302   0.6871974777902924   0.6370097776308332   0.22388227954390036   0.4841880953100143   0.08410405937797441   0.9558731978829862   0.5382204794832364   0.5918955777689546   0.012556621289219406   0.11642954743922519   0.8654698580312433   0.6986362549713458   0.554006054730737   0.4029850702325488   0.3886688980154188   0.6789496645857458   0.06895740623063015   0.26167862339078984   0.28043286175028387   0.30464206427825935
0.6389865551816762   0.47183300126894645   0.30770177393574727   0.025692421192957303   0.9517890773913839   0.8348232236381132   0.08381949439184687   0.5415043258829431   0.8676850180134095   0.8789500257551269   0.5455990149086105   0.9496087481139884   0.85512839672419   0.7625204783159018   0.6801291568773671   0.2509724931426425   0.30112234199345295   0.359535408083353   0.2914602588619483   0.5720228285568967   0.23216493576282277   0.09785678469256318   0.011027397111664434   0.2673807642786374   0.5931783805811466   0.6260237834236168   0.7033256231759172   0.24168834308568005   0.6413893031897627   0.7912005597855035   0.6195061287840703   0.700184017202737   0.7737042851763534   0.9122505340303765   0.07390711387545985   0.7505752690887486   0.9185758884521633   0.1497300557144747   0.3937779569980927   0.4996027759461061   0.6174535464587104   0.7901946476311217   0.10231769813614441   0.9275799473892093   0.38528861069588766   0.6923378629385586   0.09129030102447998   0.660199183110572   0.792110230114741   0.06631407951494185   0.3879646778485628   0.418510840024892   0.1507209269249783   0.27511351972943837   0.7684585490644925   0.718326822822155   0.377016641748625   0.3628629856990619   0.6945514351890326   0.9677515537334064   0.4584407532964616   0.21313292998458716   0.3007734781909399   0.4681487777873003
0.8409872068377512   0.4229382823534654   0.1984557800547955   0.5405688303980909   0.4556985961418636   0.7306004194149068   0.10716547903031551   0.8803696472875189   0.6635883660271226   0.664286339899965   0.7192008011817527   0.4618588072626269   0.5128674391021443   0.3891728201705267   0.9507422521172603   0.743531984440472   0.13585079735351926   0.026309834471464805   0.25619081692822765   0.7757804307070657   0.6774100440570576   0.8131769044868776   0.9554173387372877   0.3076316529197654   0.8364228372193064   0.3902386221334122   0.7569615586824923   0.7670628225216745   0.38072424107744285   0.6596382027185054   0.6497960796521767   0.8866931752341556   0.7171358750503204   0.9953518628185403   0.930595278470424   0.4248343679715287   0.20426843594817612   0.6061790426480136   0.9798530263531637   0.6813023835310567   0.06841763859465685   0.5798692081765489   0.7236622094249361   0.9055219528239911   0.3910075945375992   0.7666923036896712   0.7682448706876484   0.5978902999042256   0.5545847573182928   0.37645368155625897   0.011283312005156162   0.8308274773825511   0.17386051624084992   0.7168154788377537   0.3614872323529794   0.9441343021483956   0.4567246411905296   0.7214636160192133   0.4308919538825554   0.5192999341768668   0.25245620524235346   0.1152845733711997   0.4510389275293917   0.8379975506458102
0.1840385666476966   0.5354153651946508   0.7273767181044556   0.9324755978218191   0.7930309721100974   0.7687230615049797   0.9591318474168071   0.3345852979175935   0.2384462147918046   0.39226937994872074   0.947848535411651   0.5037578205350424   0.06458569855095471   0.6754539011109671   0.5863613030586715   0.5596235183866468   0.6078610573604252   0.9539902850917538   0.15546934917611613   0.04032358420977997   0.3554048521180717   0.8387057117205541   0.7044304216467244   0.20232603356396978   0.17136628547037508   0.3032903465259032   0.9770537035422688   0.2698504357421506   0.3783353133602777   0.5345672850209235   0.01792185612546172   0.9352651378245571   0.13988909856847306   0.14229790507220277   0.07007332071381073   0.43150731728951475   0.07530340001751837   0.46684400396123565   0.48371201765513916   0.8718837989028679   0.4674423426570932   0.512853718869482   0.32824266847902306   0.8315602146930879   0.11203749053902154   0.6741480071489279   0.6238122468322986   0.6292341811291182   0.9406712050686464   0.3708576606230246   0.6467585432900297   0.35938374538696755   0.5623358917083687   0.8362903756021011   0.628836687164568   0.42411860756241043   0.4224467931398957   0.6939924705298983   0.5587633664507573   0.9926112902728956   0.3471433931223773   0.2271484665686626   0.0750513487956181   0.12072749137002772
0.8797010504652841   0.7142947476991807   0.7468086803165951   0.28916727667693976   0.7676635599262626   0.040146740550252906   0.12299643348429648   0.6599330955478216   0.8269923548576161   0.6692890799272283   0.47623789019426677   0.30054935016085405   0.26465646314924735   0.8329987043251272   0.8474012030296988   0.8764307425984437   0.8422096700093517   0.13900623379522892   0.28863783657894154   0.883819452325548   0.4950662768869743   0.9118577672265663   0.21358648778332343   0.7630919609555202   0.6153652264216902   0.19756301952738559   0.46677780746672837   0.4739246842785805   0.8477016664954277   0.15741627897713267   0.3437813739824319   0.8139915887307589   0.02070931163781161   0.48812719904990437   0.8675434837881651   0.5134422385699048   0.7560528484885642   0.6551284947247772   0.020142280758466333   0.6370114959714612   0.9138431784792127   0.5161222609295483   0.7315044441795248   0.7531920436459132   0.41877690159223835   0.604264493702982   0.5179179563962014   0.990100082690393   0.8034116751705481   0.4067014741755964   0.051140148929473   0.5161753984118125   0.9557100086751205   0.24928519519846368   0.7073587749470411   0.7021838096810535   0.9350006970373088   0.7611579961485593   0.839815291158876   0.18874157111114873   0.17894784854874451   0.10602950142378215   0.8196730104004096   0.5517300751396875
0.26510467006953187   0.5899072404942339   0.08816856622088484   0.7985380314937743   0.8463277684772935   0.985642746791252   0.5702506098246835   0.8084379488033814   0.042916093306745416   0.5789412726156556   0.5191104608952105   0.29226255039156895   0.087206084631625   0.3296560774171919   0.8117516859481694   0.5900787407105154   0.1522053875943162   0.5684980812686325   0.9719363947892934   0.40133716959936666   0.9732575390455717   0.46246857984485046   0.15226338438888373   0.8496070944596792   0.7081528689760398   0.8725613393506165   0.06409481816799889   0.05106906296590483   0.8618251004987463   0.8869185925593646   0.49384420834331544   0.24263111416252345   0.8189090071920009   0.30797731994370897   0.9747337474481049   0.9503685637709545   0.731702922560376   0.9783212425265171   0.16298206149993558   0.3602898230604391   0.5794975349660597   0.4098231612578845   0.1910456667106422   0.9589526534610724   0.606239995920488   0.947354581413034   0.03878228232175845   0.10934555900139326   0.8980871269444481   0.07479324206241748   0.9746874641537595   0.05827649603548843   0.036262026445701825   0.1878746495030529   0.4808432558104441   0.815645381872965   0.2173530192537009   0.879897329559344   0.5061095083623391   0.8652768181020105   0.485650096693325   0.9015760870328269   0.3431274468624036   0.5049869950415714
0.9061525617272653   0.49175292577494245   0.15208178015176144   0.546034341580499   0.29991256580677733   0.5443983443619084   0.113299497830003   0.43668878257910576   0.4018254388623292   0.46960510229949093   0.13861203367624345   0.3784122865436173   0.3655634124166273   0.281730452796438   0.6577687778657993   0.5627669046706524   0.14821039316292642   0.4018331232370941   0.15165926950346012   0.6974900865686419   0.6625602964696015   0.5002570362042672   0.8085318226410565   0.1925030915270704   0.7564077347423361   0.008504110429324759   0.6564500424892951   0.6464687499465714   0.4564951689355588   0.4641057660674163   0.543150544659292   0.20977996736746565   0.05466973007322963   0.9945006637679255   0.4045385109830486   0.8313676808238484   0.6891063176566022   0.7127702109714874   0.7467697331172493   0.268600776153196   0.5408959244936759   0.3109370877343933   0.5951104636137892   0.5711106895845541   0.8783356280240744   0.8106800515301261   0.7865786409727327   0.3786075980574838   0.12192789328173832   0.8021759411008014   0.13012859848343764   0.7321388481109123   0.6654327243461795   0.33807017503338505   0.5869780538241456   0.5223588807434467   0.6107629942729499   0.3435695112654596   0.18243954284109695   0.6909911999195983   0.9216566766163476   0.6307993002939722   0.43566980972384767   0.42239042376640235
0.38076075212267174   0.3198622125595789   0.8405593461100584   0.8512797341818482   0.5024251240985973   0.5091821610294528   0.05398070513732576   0.47267213612436443   0.380497230816859   0.7070062199286514   0.9238521066538881   0.7405332880134521   0.7150645064706794   0.3689360448952663   0.33687405282974253   0.21817440727000534   0.10430151219772957   0.025366533629806728   0.15443450998864555   0.527183207350407   0.18264483558138195   0.3945672333358345   0.7187647002647979   0.10479278358400461   0.8018840834587102   0.07470502077625563   0.8782053541547394   0.2535130494021564   0.29945895936011285   0.5655228597468028   0.8242246490174137   0.780840913277792   0.9189617285432539   0.8585166398181515   0.9003725423635256   0.04030762526433997   0.2038972220725744   0.48958059492288514   0.563498489533783   0.8221332179943346   0.09959570987484484   0.4642140612930784   0.40906397954513746   0.2949500106439277   0.9169508742934629   0.0696468279572439   0.6902992792803396   0.19015722705992305   0.1150667908347527   0.9949418071809882   0.8120939251256001   0.9366441776577666   0.8156078314746398   0.4294189474341854   0.9878692761081864   0.1558032643799746   0.8966461029313859   0.5709023076160339   0.08749673374466087   0.11549563911563462   0.6927488808588116   0.08132171269314878   0.5239982442108778   0.2933624211213
0.5931531709839667   0.6171076514000704   0.11493426466574033   0.9984124104773723   0.6762022966905038   0.5474608234428264   0.42463498538540073   0.8082551834174493   0.5611355058557511   0.5525190162618382   0.6125410602598006   0.8716110057596826   0.7455276743811113   0.12310006882765274   0.6246717841516142   0.715807741379708   0.8488815714497253   0.5521977612116188   0.5371750504069533   0.6003121022640734   0.15613269059091378   0.47087604851847004   0.013176806196075499   0.30694968114277343   0.562979519606947   0.8537683971183997   0.8982425415303351   0.3085372706654011   0.8867772229164432   0.3063075736755732   0.4736075561449344   0.5002820872479518   0.3256417170606921   0.7537885574137351   0.8610664958851337   0.6286710814882692   0.5801140426795808   0.6306884885860823   0.23639471173351959   0.9128633401085612   0.7312324712298555   0.07849072737446351   0.6992196613265663   0.31255123784448774   0.5750997806389417   0.6076146788559935   0.6860428551304908   0.005601556701714331   0.012120261031994645   0.7538462817375938   0.7878003136001556   0.6970642860363132   0.12534303811555142   0.44753870806202056   0.3141927574552212   0.19678219878836145   0.7997013210548594   0.6937501506482855   0.45312626157008745   0.5681111173000922   0.2195872783752785   0.06306166206220316   0.21673154983656784   0.6552477771915312
0.488354807145423   0.9845709346877396   0.5175118885100015   0.3426965393470434   0.9132550265064813   0.3769562558317462   0.8314690333795108   0.33709498264532906   0.9011347654744867   0.6231099740941524   0.043668719779355165   0.6400306966090158   0.7757917273589353   0.1755712660321318   0.7294759623241339   0.44324849782065434   0.976090406304076   0.4818211153838463   0.2763497007540465   0.8751373805205621   0.7565031279287975   0.4187594533216431   0.059618150917478706   0.21988960332903096   0.2681483207833744   0.43418851863390345   0.5421062624074772   0.8771930639819876   0.3548932942768931   0.057232262802157305   0.7106372290279663   0.5400980813366585   0.4537585288024064   0.43412228870800496   0.6669685092486112   0.9000673847276427   0.6779668014434712   0.25855102267587315   0.9374925469244773   0.45681888690698835   0.7018763951393953   0.7767299072920268   0.6611428461704307   0.5816815063864262   0.9453732672105978   0.35797045397038374   0.601524695252952   0.3617919030573953   0.6772249464272233   0.9237819353364802   0.05941843284547484   0.4845988390754077   0.3223316521503302   0.8665496725343229   0.3487812038175085   0.9445007577387492   0.8685731233479238   0.432427383826318   0.6818126945688973   0.044433373011106454   0.19060632190445262   0.17387636115044489   0.74432014764442   0.5876144861041181
0.4887299267650574   0.397146453858418   0.08317730147398934   0.005932979717691852   0.5433566595544597   0.0391759998880343   0.48165260622103734   0.6441410766602965   0.8661317131272362   0.11539406455155404   0.4222341733755625   0.15954223758488886   0.543800060976906   0.2488443920172311   0.07345296955805403   0.2150414798461397   0.6752269376289822   0.8164170081909131   0.39164027498915677   0.17060810683503325   0.48462061572452964   0.6425406470404682   0.6473201273447368   0.5829936207309151   0.9958906889594723   0.2453941931820502   0.5641428258707474   0.5770606410132233   0.45253402940501264   0.2062181932940159   0.08249021964971003   0.9329195643529267   0.5864023162777764   0.09082412874246183   0.6602560462741475   0.7733773267680378   0.04260225530087032   0.8419797367252307   0.5868030767160934   0.5583358469218982   0.367375317671888   0.025562728534317663   0.19516280172693673   0.3877277400868649   0.8827547019473584   0.3830220814938495   0.5478426743822   0.8047341193559497   0.8868640129878861   0.13762788831179928   0.9836998485114526   0.22767347834272647   0.43432998358287345   0.9314096950177834   0.9012096288617426   0.2947539139897998   0.847927667305097   0.8405855662753215   0.2409535825875951   0.521376587221762   0.8053254120042268   0.9986058295500908   0.6541505058715016   0.9630407402998638
0.4379500943323387   0.9730431010157732   0.4589877041445649   0.5753130002129989   0.5551953923849803   0.5900210195219237   0.9111450297623649   0.7705788808570491   0.6683313793970942   0.4523931312101244   0.9274451812509122   0.5429054025143226   0.23400139581422078   0.520983436192341   0.026235552389169615   0.24815148852452287   0.3860737285091237   0.6803978699170194   0.7852819698015745   0.7267749013027609   0.5807483165048969   0.6817920403669286   0.13113146393007286   0.7637341610028971   0.14279822217255822   0.7087489393511555   0.672143759785508   0.18842116078989832   0.5876028297875779   0.11872791982923177   0.7609987300231431   0.4178422799328492   0.9192714503904837   0.6663347886191073   0.8335535487722309   0.8749368774185265   0.6852700545762629   0.14535135242676633   0.8073179963830612   0.6267853888940037   0.29919632606713925   0.4649534825097469   0.02203602658148672   0.9000104875912428   0.7184480095622423   0.7831614421428182   0.8909045626514138   0.1362763265883456   0.5756497873896841   0.07441250279166275   0.21876080286590588   0.9478551657984473   0.9880469576021061   0.955684582962431   0.4577620728427628   0.530012885865598   0.06877550721162247   0.28934979434332364   0.624208524070532   0.6550760084470715   0.3835054526353595   0.14399844191655733   0.8168905276874707   0.02829061955306774
0.08430912656822029   0.6790449594068104   0.794854501105984   0.12828013196182494   0.365861117005978   0.8958835172639922   0.9039499384545702   0.9920038053734793   0.7902113296162939   0.8214710144723295   0.6851891355886643   0.044148639575032046   0.8021643720141878   0.8657864315098984   0.22742706274590146   0.514135753709434   0.7333888648025653   0.5764366371665748   0.6032185386753695   0.8590597452623625   0.34988341216720575   0.43243819525001753   0.7863280109878987   0.8307691257092947   0.26557428559898544   0.753393235843207   0.9914735098819147   0.7024889937474698   0.8997131685930074   0.8575097185792149   0.08752357142734452   0.7104851883739904   0.10950183897671356   0.03603870410688536   0.4023344358386802   0.6663365487989584   0.3073374669625258   0.1702522725969869   0.17490737309277873   0.15220079508952444   0.5739486021599606   0.593815635430412   0.5716888344174093   0.29314104982716194   0.22406518999275477   0.16137744018039454   0.7853608234295105   0.4623719241178672   0.9584909043937693   0.40798420433718746   0.7938873135475958   0.7598829303703973   0.05877773580076184   0.5504744857579726   0.7063637421202513   0.04939774199640692   0.9492758968240483   0.5144357816510873   0.3040293062815711   0.3830611931974485   0.6419384298615225   0.3441835090541004   0.12912193318879234   0.23086039810792405
0.06798982770156195   0.7503678736236884   0.5574330987713831   0.9377193482807621   0.8439246377088072   0.5889904334432938   0.7720722753418726   0.4753474241628949   0.8854337333150378   0.18100622910610634   0.9781849617942768   0.7154644937924975   0.826655997514276   0.6305317433481337   0.2718212196740255   0.6660667517960907   0.8773801006902278   0.11609596169704639   0.9677919133924544   0.2830055585986421   0.23544167082870526   0.771912452642946   0.838669980203662   0.05214516049071806   0.1674518431271433   0.02154457901925761   0.281236881432279   0.11442581220995596   0.32352720541833613   0.4325541455759638   0.5091646060904064   0.6390783880470611   0.4380934721032983   0.2515479164698574   0.5309796442961296   0.9236138942545635   0.6114374745890223   0.6210161731217237   0.2591584246221041   0.25754714245847293   0.7340573738987946   0.5049202114246774   0.2913665112296497   0.9745415838598308   0.4986157030700893   0.7330077587817314   0.45269653102598767   0.9223964233691128   0.33116385994294595   0.7114631797624738   0.17145964959370869   0.8079706111591568   0.007636654524609831   0.27890903418651   0.6622950435033023   0.16889222311209576   0.5695431824213115   0.027361117716652547   0.1313153992071727   0.2452783288575322   0.9581057078322893   0.4063449445949288   0.8721569745850686   0.9877311863990593
0.22404833393349474   0.9014247331702514   0.5807904633554188   0.01318960253922847   0.7254326308634055   0.16841697438852007   0.12809393232943123   0.09079317917011571   0.3942687709204595   0.4569537946260463   0.9566342827357226   0.2828225680109589   0.38663211639584966   0.17804476043953632   0.2943392392324203   0.11393034489886317   0.8170889339745381   0.15068364272288376   0.16302384002524756   0.8686520160413309   0.8589832261422489   0.744338698127955   0.290866865440179   0.8809208296422717   0.6349348922087541   0.8429139649577035   0.7100764020847601   0.8677312271030432   0.9095022613453486   0.6744969905691834   0.5819824697553289   0.7769380479329275   0.5152334904248891   0.21754319594313715   0.6253481870196063   0.4941154799219686   0.12860137402903946   0.03949843550360084   0.33100894778718604   0.3801851350231054   0.31151244005450135   0.8888147927807171   0.1679851077619385   0.5115331189817744   0.4525292139122525   0.1444760946527621   0.8771182423217595   0.6306122893395028   0.8175943217034984   0.3015621296950586   0.16704184023699944   0.7628810622364596   0.9080920603581498   0.6270651391258751   0.5850593704816706   0.985943014303532   0.3928585699332607   0.409521943182738   0.9597111834620643   0.4918275343815635   0.2642571959042212   0.3700235076791371   0.6287022356748782   0.11164239935845811
0.9527447558497198   0.48120871489842004   0.4607171279129397   0.6001092803766837   0.5002155419374673   0.336732620245658   0.5835988855911801   0.9694969910371809   0.682621220233969   0.035170490550599384   0.4165570453541807   0.20661592880072133   0.7745291598758192   0.40810535142472426   0.8314976748725101   0.22067291449718926   0.3816705899425585   0.9985834082419863   0.8717864914104458   0.7288453801156257   0.11741339403833728   0.6285599005628492   0.2430842557355677   0.6172029807571676   0.16466863818861743   0.1473511856644291   0.782367127822628   0.017093700380483936   0.6644530962511501   0.8106185654187711   0.19876824223144782   0.047596709343303026   0.9818318760171811   0.7754480748681717   0.7822111968772671   0.8409807805425817   0.20730271614136198   0.3673427234434475   0.9507135220047569   0.6203078660453925   0.8256321261988034   0.3687593152014612   0.07892703059431105   0.8914624859297667   0.7082187321604662   0.740199414638612   0.8358427748587434   0.2742595051725991   0.5435500939718487   0.592848228974183   0.05347564703611539   0.25716580479211515   0.8790969977206987   0.7822296635554118   0.8547074048046676   0.20956909544881214   0.8972651217035176   0.006781588687240083   0.07249620792740047   0.36858831490623045   0.6899624055621556   0.6394388652437926   0.12178268592264353   0.748280448860838
0.8643302793633522   0.2706795500423314   0.04285565532833248   0.8568179629310713   0.15611154720288595   0.5304801354037194   0.2070128804695891   0.5825584577584721   0.6125614532310372   0.9376319064295364   0.15353723343347372   0.325392652966357   0.7334644555103386   0.1554022428741246   0.29882982862880614   0.11582355751754488   0.836199333806821   0.14862065418688453   0.22633362070140567   0.7472352426113145   0.14623692824466533   0.509181788943092   0.10455093477876215   0.9989547937504765   0.2819066488813132   0.2385022389007605   0.06169527945042967   0.14213683081940515   0.12579510167842725   0.7080221034970411   0.8546823989808405   0.5595783730609329   0.5132336484473901   0.7703901970675047   0.7011451655473668   0.23418572009457594   0.7797691929370515   0.61498795419338   0.4023153369185607   0.11836216257703108   0.9435698591302306   0.46636730000649557   0.17598171621715503   0.3711269199657167   0.7973329308855652   0.9571855110634037   0.07143078143839288   0.3721721262152402   0.5154262820042521   0.7186832721626432   0.009735501987963203   0.2300352953958351   0.38963118032582483   0.010661168665601985   0.15505310300712263   0.6704569223349022   0.8763975318784347   0.2402709715980973   0.4539079374597558   0.4362712022403262   0.09662833894138323   0.6252830174047173   0.05159260054119509   0.3179090396632951
0.15305847981115264   0.15891571739822166   0.8756108843240401   0.9467821196975784   0.3557255489255874   0.20173020633481806   0.8041801028856472   0.5746099934823382   0.8402992669213353   0.4830469341721749   0.794444600897684   0.34457469808650315   0.4506680865955105   0.47238576550657296   0.6393914978905614   0.674117775751601   0.5742705547170758   0.23211479390847567   0.18548356043080558   0.23784657351127483   0.4776422157756925   0.6068317765037584   0.13389095988961047   0.9199375338479797   0.3245837359645399   0.4479160591055368   0.2582800755655704   0.9731554141504013   0.9688581870389524   0.24618585277071872   0.4540999726799232   0.3985454206680631   0.12855892011761716   0.7631389185985438   0.6596553717822392   0.05397072258155993   0.6778908335221067   0.2907531530919708   0.02026387389167785   0.3798529468299589   0.10362027880503091   0.05863835918349515   0.8347803134608723   0.14200637331868407   0.6259780630293384   0.4518065826797367   0.7008893535712618   0.22206883947070433   0.3013943270647985   0.003890523574199936   0.4426092780056914   0.24891342532030303   0.3325361400258461   0.7577046708034813   0.9885093053257682   0.8503680046522399   0.2039772199082289   0.9945657522049375   0.328853933543529   0.7963972820706801   0.5260863863861223   0.7038125991129667   0.30859005965185116   0.4165443352407211
0.4224661075810914   0.6451742399294714   0.4738097461909789   0.27453796192203705   0.7964880445517529   0.19336765724973476   0.772920392619717   0.05246912245133273   0.4950937174869544   0.18947713367553481   0.3303111146140256   0.8035556971310297   0.16255757746110835   0.4317724628720536   0.34180180928825743   0.9531876924787898   0.9585803575528794   0.4372067106671162   0.012947875744728447   0.1567904104081097   0.4324939711667572   0.7333941115541496   0.7043578160928773   0.7402460751673886   0.01002786358566584   0.08821987162467806   0.23054806990189844   0.4657081132453515   0.2135398190339129   0.8948522143749433   0.4576276772821814   0.41323899079401877   0.7184461015469585   0.7053750806994085   0.12731656266815575   0.6096832936629891   0.5558885240858501   0.27360261782735484   0.7855147533798983   0.6564956011841994   0.5973081665329707   0.8363959071602387   0.7725668776351698   0.49970519077608966   0.1648141953662135   0.10300179560608916   0.06820906154229255   0.759459115608701   0.15478633178054765   0.014781923981411088   0.8376609916403941   0.29375100236334956   0.9412465127466347   0.11992970960646779   0.38003331435821275   0.8805120115693308   0.22280041119967628   0.4145546289070593   0.252716751690057   0.27082871790634166   0.6669118871138261   0.14095201107970445   0.4672019983101587   0.6143331167221423
0.06960372058085545   0.30455610391946575   0.6946351206749888   0.11462792594605266   0.904789525214642   0.2015543083133766   0.6264260591326962   0.3551688103373516   0.7500031934340943   0.1867723843319655   0.7887650674923021   0.061417807974002   0.8087566806874595   0.06684267472549772   0.40873175313408944   0.18090579640467122   0.5859562694877832   0.6522880458184384   0.15601500144403246   0.9100770784983295   0.9190443823739571   0.511336034738734   0.6888130031338738   0.2957439617761872   0.8494406617931016   0.2067799308192682   0.9941778824588849   0.18111603583013455   0.9446511365784597   0.005225622505891624   0.36775182332618866   0.825947225492783   0.1946479431443654   0.8184532381739261   0.5789867558338865   0.764529417518781   0.3858912624569058   0.7516105634484284   0.17025500269979707   0.5836236211141097   0.7999349929691225   0.09932251762998999   0.0142400012557646   0.6735465426157802   0.8808906105951654   0.587986482891256   0.3254269981218908   0.377802580839593   0.031449948802063754   0.38120655207198784   0.33124911566300586   0.19668654500945845   0.08679881222360405   0.3759809295660962   0.9634972923368171   0.3707393195166755   0.8921508690792387   0.5575276913921701   0.38451053650293066   0.6062099019978945   0.5062596066223328   0.8059171279437417   0.21425553380313359   0.02258628088378477
0.7063246136532103   0.7065946103137517   0.200015532547369   0.34903973826800455   0.8254340030580448   0.11860812742249564   0.8745885344254781   0.9712371574284115   0.7939840542559811   0.7374015753505079   0.5433394187624723   0.7745506124189531   0.7071852420323771   0.36142064578441163   0.5798421264256551   0.40381129290227763   0.8150343729531384   0.8038929543922415   0.19533158992272448   0.7976013909043831   0.30877476633080553   0.9979758264484999   0.9810760561195909   0.7750151100205983   0.6024501526775953   0.2913812161347482   0.7810605235722219   0.4259753717525938   0.7770161496195503   0.17277308871225258   0.9064719891467438   0.4547382143241822   0.9830320953635693   0.43537151336174473   0.3631325703842714   0.6801876019052291   0.27584685333119224   0.07395086757733312   0.7832904439586162   0.27637630900295146   0.46081248037805383   0.27005791318509154   0.5879588540358918   0.4787749180985683   0.15203771404724833   0.2720820867365917   0.6068827979163008   0.70375980807797   0.549587561369653   0.9807008706018434   0.825822274344079   0.2777844363253762   0.7725714117501027   0.8079277818895909   0.9193502851973353   0.8230462220011939   0.7895393163865334   0.3725562685278461   0.5562177148130639   0.1428586200959649   0.5136924630553411   0.298605400950513   0.7729272708544477   0.8664823110930134
0.0528799826772873   0.028547487765421452   0.1849684168185559   0.38770739299444507   0.900842268630039   0.7564654010288298   0.578085618902255   0.6839475849164751   0.35125470726038593   0.7757645304269863   0.752263344558176   0.4061631485910989   0.5786832955102832   0.9678367485373955   0.8329130593608407   0.5831169265899049   0.7891439791237498   0.5952804800095494   0.2766953445477769   0.44025830649394004   0.2754515160684087   0.2966750790590364   0.5037680736933292   0.5737759954009266   0.22257153339112137   0.2681275912936149   0.31879965687477335   0.18606860240648151   0.3217292647610824   0.5116621902647851   0.7407140379725183   0.5021210174900065   0.9704745575006964   0.7358976598377988   0.9884506934143423   0.09595786889890753   0.39179126199041325   0.7680609113004033   0.15553763405350154   0.5128409423090027   0.6026472828666634   0.1727804312908539   0.8788422895057247   0.0725826358150626   0.32719576679825474   0.8761053522318175   0.3750742158123955   0.49880664041413597   0.10462423340713337   0.6079777609382025   0.056274558937622114   0.3127380380076545   0.782894968646051   0.09631557067341746   0.3155605209651038   0.8106170205176481   0.8124204111453545   0.3604179108356187   0.32710982755076146   0.7146591516187405   0.42062914915494126   0.5923569995352154   0.1715721934972599   0.20181820930973787
0.8179818662882778   0.4195765682443615   0.2927299039915352   0.12923557349467527   0.4907860994900231   0.543471216012544   0.9176556881791398   0.6304289330805393   0.3861618660828897   0.9354934550743413   0.8613811292415177   0.31769089507288484   0.6032668974368387   0.8391778844009239   0.5458206082764139   0.5070738745552368   0.7908464862914842   0.4787599735653052   0.2187107807256524   0.7924147229364963   0.370217337136543   0.8864029740300898   0.04713858722839249   0.5905965136267585   0.5522354708482652   0.4668264057857283   0.7544086832368573   0.4613609401320832   0.06144937135824207   0.9233551897731844   0.8367529950577175   0.8309320070515439   0.6752875052753523   0.987861734698843   0.9753718658161998   0.5132411119786591   0.07202060783851359   0.1486838502979191   0.42955125753978596   0.0061672374234222685   0.2811741215470293   0.6699238767326139   0.21084047681413357   0.21375251448692598   0.9109567844104863   0.7835209027025241   0.16370188958574108   0.6231560008601675   0.35872131356222114   0.31669449691679574   0.40929320634888383   0.16179506072808436   0.29727194220397907   0.3933393071436113   0.5725402112911663   0.3308630536765405   0.6219844369286267   0.40547757244476834   0.5971683454749664   0.8176219416978814   0.5499638290901132   0.2567937221468492   0.16761708793518051   0.8114547042744592
0.26878970754308384   0.5868698454142354   0.956776611121047   0.5977021897875332   0.3578329231325975   0.8033489427117113   0.7930747215353059   0.9745461889273657   0.9991116095703764   0.48665444579491557   0.38378151518642206   0.8127511281992813   0.7018396673663972   0.09331513865130422   0.8112413038952557   0.4818880745227408   0.07985523043777049   0.6878375662065359   0.21407295842028928   0.6642661328248594   0.5298914013476573   0.43104384405968665   0.04645587048510876   0.8528114285504002   0.2611016938045735   0.8441739986454513   0.0896792593640618   0.255109238762867   0.903268770671976   0.04082505593374005   0.2966045378287559   0.28056304983550134   0.9041571611015997   0.5541706101388245   0.9128230226423338   0.46781192163622004   0.2023174937352024   0.46085547148752026   0.1015817187470781   0.9859238471134792   0.12246226329743193   0.7730179052809844   0.8875087603267888   0.3216577142886199   0.5925708619497746   0.3419740612212977   0.84105288984168   0.46884628573821974   0.3314691681452011   0.49780006257584636   0.7513736304776183   0.21373704697535273   0.4282003974732251   0.45697500664210633   0.45476909264886234   0.9331739971398514   0.5240432363716254   0.9028043965032818   0.5419460700065285   0.46536207550363134   0.321725742636423   0.44194892501576155   0.4403643512594504   0.4794382283901521
0.19926347933899108   0.6689310197347772   0.5528555909326616   0.15778051410153218   0.6066926173892164   0.3269569585134795   0.7118027010909815   0.6889342283633124   0.2752234492440154   0.8291568959376331   0.9604290706133632   0.47519718138795974   0.8470230517707903   0.3721818892955268   0.5056599779645009   0.5420231842481084   0.32297981539916487   0.46937749279224494   0.9637139079579725   0.07666110874447701   0.0012540727627418393   0.027428567776483403   0.5233495566985221   0.5972228803543249   0.8019905934237508   0.3584975480417062   0.9704939657658606   0.43944236625279276   0.1952979760345343   0.03154058952822671   0.258691264674879   0.7505081378894802   0.9200745267905189   0.2023836935905936   0.2982621940615158   0.27531095650152054   0.07305147501972864   0.8302018042950668   0.7926022160970149   0.7332877722534121   0.7500716596205638   0.36082431150282185   0.8288883081390424   0.6566266635089352   0.748817586857822   0.3333957437263384   0.30553875144052023   0.059403783154610236   0.9468269934340712   0.9748981956846322   0.33504478567465973   0.6199614169018175   0.7515290173995369   0.9433576061564055   0.07635352099978068   0.8694532790123373   0.831454490609018   0.7409739125658119   0.7780913269382649   0.5941423225108167   0.7584030155892894   0.9107721082707451   0.9854891108412501   0.8608545502574045
0.008331355968725545   0.5499477967679233   0.15660080270220772   0.2042278867484694   0.25951376911090357   0.21655205304158487   0.8510620512616874   0.14482410359385917   0.3126867756768324   0.24165385735695266   0.5160172655870278   0.5248626866920416   0.5611577582772955   0.29829625120054715   0.4396637445872471   0.6554094076797045   0.7297032676682775   0.5573223386347352   0.6615724176489822   0.06126708516888771   0.9713002520789882   0.6465502303639902   0.6760833068077321   0.20041253491148317   0.9629688961102626   0.09660243359606685   0.5194825041055243   0.9961846481630138   0.7034551269993591   0.8800503805544819   0.6684204528438369   0.8513605445691546   0.39076835132252663   0.6383965231975294   0.15240318725680913   0.32649785787711294   0.8296105930452311   0.3401002719969822   0.712739442669562   0.6710884501974085   0.09990732537695364   0.7827779333622469   0.051167025020579855   0.6098213650285208   0.12860707329796547   0.1362277029982568   0.37508371821284775   0.40940883011703766   0.16563817718770285   0.03962526940218994   0.8556012141073234   0.4132241819540239   0.4621830501883438   0.15957488884770796   0.18718076126348648   0.5618636373848693   0.07141469886581718   0.5211783656501786   0.03477757400667736   0.23536577950775633   0.24180410582058603   0.18107809365319646   0.32203813133711534   0.5642773293103478
0.14189678044363238   0.39830016029094956   0.27087110631653544   0.954455964281827   0.013289707145666919   0.26207245729269274   0.8957873881036877   0.5450471341647893   0.8476515299579641   0.22244718789050283   0.04018617399636432   0.13182295221076545   0.38546847976962023   0.06287229904279486   0.8530054127328779   0.5699593148258961   0.3140537809038031   0.5416939333926162   0.8182278387262005   0.3345935353181398   0.07224967508321703   0.36061583973941974   0.4961897073890852   0.7703162060077919   0.9303528946395846   0.9623156794484702   0.2253186010725497   0.8158602417259649   0.9170631874939177   0.7002432221557774   0.329531212968862   0.27081310756117566   0.06941165753595366   0.4777960342652746   0.2893450389724977   0.13899015535041018   0.6839431777663334   0.4149237352224798   0.4363396262396198   0.569030840524514   0.36988939686253036   0.8732298018298635   0.6181117875134193   0.2344373052063742   0.2976397217793133   0.5126139620904439   0.12192208012433418   0.46412109919858224   0.36728682713972866   0.5502982826419736   0.8966034790517845   0.6482608574726172   0.45022363964581097   0.8500550604861962   0.5670722660829225   0.3774477499114416   0.3808119821098573   0.37225902622092155   0.2777272271104248   0.2384575945610314   0.6968688043435239   0.9573352909984417   0.841387600870805   0.6694267540365174
0.3269794074809936   0.08410548916857821   0.22327581335738564   0.4349894488301432   0.029339685701680246   0.5714915270781344   0.10135373323305144   0.970868349631561   0.6620528585619516   0.021193244436160812   0.20475025418126697   0.3226074921589437   0.21182921891614062   0.17113818394996466   0.6376779880983445   0.9451597422475021   0.8310172368062834   0.7988791577290432   0.35995076098791967   0.7067021476864707   0.13414843246275943   0.8415438667306013   0.5185631601171147   0.037275393649953296   0.8071690249817659   0.7574383775620231   0.29528734675972906   0.6022859448198101   0.7778293392800856   0.18594685048388873   0.19393361352667762   0.6314175951882491   0.11577648071813404   0.16475360604772793   0.9891833593454107   0.30881010302930545   0.9039472618019935   0.9936154220977633   0.35150537124706616   0.36365036078180335   0.0729300249957101   0.19473626436872016   0.9915546102591465   0.6569482130953327   0.9387815925329507   0.35319239763811877   0.47299145014203176   0.6196728194453793   0.1316125675511848   0.5957540200760957   0.1777041033823027   0.01738687462556923   0.3537832282710992   0.40980716959220687   0.9837704898556251   0.38596927943732007   0.23800674755296516   0.24505356354447896   0.9945871305102144   0.07715917640801462   0.3340594857509717   0.25143814144671567   0.6430817592631483   0.7135088156262113
0.26112946075526167   0.056701877077995545   0.6515271490040018   0.05656060253087863   0.322347868222311   0.7035094794398767   0.17853569886196996   0.4368877830854993   0.19073530067112615   0.10775545936378113   0.0008315954796672788   0.41950090845993004   0.8369520724000269   0.6979482897715742   0.01706110562404222   0.03353162902260999   0.5989453248470618   0.45289472622709526   0.022473975113827826   0.9563724526145954   0.26488583909609004   0.2014565847803796   0.3793922158506796   0.2428636369883841   0.003756378340828399   0.14475470770238405   0.7278650668466778   0.18630303445750546   0.6814085101185174   0.4412452282625073   0.5493293679847079   0.7494152513720062   0.4906732094473913   0.33348976889872617   0.5484977725050406   0.3299143429120761   0.6537211370473643   0.6355414791271519   0.5314366668809983   0.29638271388946613   0.054775812200302566   0.18264675290005664   0.5089626917671706   0.3400102612748708   0.7898899731042125   0.9811901681196771   0.12957047591649096   0.09714662428648668   0.7861335947633842   0.836435460417293   0.4017054090698131   0.9108435898289812   0.10472508464486668   0.3951902321547857   0.8523760410851052   0.16142833845697502   0.6140518751974754   0.06170046325605956   0.3038782685800646   0.8315139955448989   0.960330738150111   0.4261589841289077   0.7724416016990662   0.5351312816554328
0.9055549259498085   0.24351223122885102   0.26347890993189566   0.19512102038056198   0.11566495284559596   0.262322063109174   0.1339084340154047   0.09797439609407528   0.32953135808221184   0.425886602691881   0.7322030249455916   0.18713080626509407   0.22480627343734513   0.030696370537095292   0.8798269838604864   0.02570246780811905   0.6107543982398698   0.9689959072810357   0.5759487152804218   0.19418847226322017   0.6504236600897587   0.5428369231521281   0.8035071135813555   0.6590571906077874   0.7448687341399503   0.29932469192327704   0.5400282036494599   0.46393617022722544   0.6292037812943543   0.03700262881410306   0.40611976963405516   0.3659617741331502   0.29967242321214244   0.611116026122222   0.6739167446884636   0.1788309678680561   0.07486614977479729   0.5804196555851268   0.7940897608279772   0.15312850005993706   0.46411175153492756   0.6114237483040911   0.21814104554755542   0.9589400277967168   0.8136880914451688   0.06858682515196295   0.4146339319661999   0.29988283718892944   0.06881935730521863   0.7692621332286859   0.87460572831674   0.8359466669617039   0.4396155760108644   0.7322595044145829   0.46848595868268483   0.4699848928285538   0.13994315279872194   0.12114347829236079   0.7945692139942212   0.29115392496049775   0.06507700302392465   0.5407238227072341   0.00047945316624402714   0.1380254249005607
0.6009652514889972   0.929300074403143   0.7823384076186886   0.1790853971038438   0.7872771600438283   0.8607132492511801   0.3677044756524887   0.8792025599149144   0.7184578027386096   0.09145111602249414   0.4930987473357487   0.043255892953210355   0.2788422267277453   0.3591916116079113   0.024612788653063895   0.5732710001246565   0.13889907392902334   0.23804813331555053   0.23004357465884268   0.2821170751641588   0.07382207090509871   0.6973243106083165   0.22956412149259864   0.1440916502635981   0.4728568194161016   0.7680242362051735   0.44722571387391   0.9650062531597543   0.6855796593722734   0.9073109869539935   0.07952123822142133   0.08580369324483994   0.9671218566336637   0.8158598709314993   0.5864224908856727   0.04254780029162959   0.6882796299059184   0.456668259323588   0.5618097022326087   0.46927680016697304   0.5493805559768951   0.21862012600803746   0.33176612757376606   0.18715972500281428   0.4755584850717964   0.5212958153997209   0.10220200608116743   0.043068074739216165   0.002701665655694753   0.7532715791945475   0.6549762922072574   0.07806182157946187   0.3171220062834214   0.845960592240554   0.5754550539858361   0.9922581283346219   0.35000014964975773   0.030100721309054695   0.9890325631001634   0.9497103280429924   0.6617205197438393   0.5734324619854667   0.42722286086755473   0.4804335278760193
0.11233996376694422   0.3548123359774292   0.09545673329378865   0.293273802873205   0.6367814786951479   0.8335165205777083   0.9932547272126212   0.25020572813398884   0.6340798130394532   0.08024494138316081   0.3382784350053638   0.17214390655452697   0.3169578067560317   0.23428434914260682   0.7628233810195277   0.17988577821990503   0.966957657106274   0.20418362783355212   0.7737908179193643   0.2301754501769127   0.3052371373624347   0.6307511658480854   0.34656795705180965   0.7497419223008934   0.1928971735954905   0.2759388298706562   0.251111223758021   0.45646811942768845   0.5561156949003426   0.4424223092929479   0.25785649654539977   0.2062623912936996   0.9220358818608896   0.3621773679097871   0.919578061540036   0.034118484739172644   0.6050780751048579   0.1278930187671803   0.15675468052050817   0.8542327065192676   0.6381204179985839   0.9237093909336281   0.38296386260114385   0.6240572563423549   0.33288328063614914   0.29295822508554276   0.0363959055493342   0.8743153340414614   0.13998610704065867   0.01701939521488658   0.7852846817913132   0.417847214613773   0.583870412140316   0.5745970859219387   0.5274281852459135   0.21158482332007342   0.6618345302794265   0.21241971801215156   0.6078501237058775   0.17746633858090077   0.05675645517456865   0.08452669924497126   0.4510954431853693   0.32323363206163314
0.4186360371759848   0.16081730831134308   0.06813158058422551   0.6991763757192783   0.08575275653983563   0.8678590832258003   0.03173567503489131   0.8248610416778168   0.945766649499177   0.8508396880109137   0.24645099324357808   0.40701382706404376   0.36189623735886095   0.27624260208897505   0.7190228079976646   0.19542900374397038   0.7000617070794345   0.0638228840768235   0.11117268429178713   0.01796266516306963   0.6433052519048658   0.9792961848318522   0.6600772411064177   0.6947290331014365   0.22466921472888102   0.8184788765205092   0.5919456605221923   0.9955526573821583   0.13891645818904538   0.9506197932947089   0.5602099854873009   0.1706916157043414   0.19314980868986842   0.09978010528379513   0.3137589922437229   0.7636777886402976   0.8312535713310075   0.8235375031948201   0.5947361842460582   0.5682487848963272   0.13119186425157303   0.7597146191179965   0.4835634999542711   0.5502861197332576   0.4878866123467072   0.7804184342861443   0.8234862588478533   0.8555570866318212   0.26321739761782625   0.9619395577656351   0.23154059832566104   0.8600044292496629   0.12430093942878086   0.011319764470926273   0.67133061283836   0.6893128135453215   0.9311511307389124   0.9115396591871311   0.3575716205946372   0.9256350249050239   0.09989755940790496   0.08800215599231108   0.762835436348579   0.3573862400086967
0.9687056951563319   0.3282875368743145   0.27927193639430786   0.8071001202754391   0.4808190828096247   0.5478691025881702   0.45578567754645455   0.9515430336436179   0.21760168519179846   0.5859295448225351   0.22424507922079348   0.09153860439395503   0.09330074576301761   0.5746097803516088   0.5529144663824334   0.4022257908486335   0.16214961502410516   0.6630701211644777   0.1953428457877962   0.47659076594360966   0.06225205561620021   0.5750679651721666   0.4325074094392172   0.11920452593491297   0.09354636045986828   0.24678042829785207   0.15323547304490936   0.3121044056594739   0.6127272776502436   0.6989113257096818   0.6974497954984549   0.3605613720158559   0.39512559245844514   0.11298178088714675   0.47320471627766136   0.2690227676219009   0.30182484669542753   0.5383720005355379   0.920290249895228   0.8667969767732674   0.13967523167132237   0.8753018793710603   0.7249474041074317   0.39020621082965773   0.07742317605512215   0.30023391419889367   0.2924399946682145   0.2710016848947448   0.9838768155952539   0.053453485901041625   0.13920452162330516   0.9588972792352709   0.37114953794501027   0.3545421601913598   0.4417547261248503   0.598335907219415   0.9760239454865651   0.24156037930421304   0.968550009847189   0.329313139597514   0.6741990987911376   0.7031883787686751   0.04825975995196098   0.4625161628242466
0.5345238671198153   0.8278864993976148   0.3233123558445292   0.0723099519945889   0.4571006910646931   0.5276525851987212   0.030872361176314686   0.8013082670998442   0.4732238754694392   0.4741990992976795   0.8916678395530095   0.8424109878645732   0.10207433752442893   0.1196569391063197   0.4499131134281592   0.2440750806451583   0.12605039203786378   0.8780965598021067   0.4813631035809703   0.9147619410476443   0.4518512932467262   0.1749081810334316   0.4331033436290093   0.4522457782233976   0.917327426126911   0.34702168163581676   0.1097909877844801   0.3799358262288087   0.4602267350622179   0.8193690964370957   0.07891862660816541   0.5786275591289646   0.9870028595927787   0.34516999713941615   0.18725078705515588   0.7362165712643913   0.8849285220683497   0.22551305803309646   0.7373376736269966   0.49214149061923307   0.758878130030486   0.34741649823098975   0.25597457004602636   0.5773795495715888   0.30702683678375975   0.1725083171975582   0.822871226417017   0.1251337713481912   0.3896994106568488   0.8254866355617414   0.713080238632537   0.7451979451193825   0.929472675594631   0.0061175391246457225   0.6341616120243715   0.1665703859904179   0.9424698160018523   0.6609475419852295   0.4469108249692157   0.4303538147260265   0.05754129393350252   0.4354344839521331   0.709573151342219   0.9382123241067934
0.29866316390301656   0.08801798572114333   0.4535985812961927   0.3608327745352047   0.9916363271192568   0.9155096685235852   0.6307273548791756   0.23569900318701345   0.601936916462408   0.09002303296184377   0.9176471162466386   0.49050105806763095   0.672464240867777   0.08390549383719804   0.28348550422226715   0.32393067207721304   0.7299944248659248   0.4229579518519685   0.8365746792530514   0.8935768573511865   0.6724531309324223   0.9875234678998354   0.12700152791083244   0.9553645332443931   0.3737899670294057   0.8995054821786921   0.6734029466146397   0.5945317587091884   0.3821536399101489   0.9839958136551069   0.04267559173546415   0.3588327555221749   0.780216723447741   0.8939727806932631   0.12502847548882548   0.868331697454544   0.10775248257996387   0.8100672868560651   0.8415429712665583   0.5444010253773309   0.3777580577140391   0.3871093350040966   0.0049682920135069   0.6508241680261444   0.7053049267816168   0.3995858671042612   0.8779667641026745   0.6954596347817513   0.33151495975221107   0.5000803849255692   0.2045638174880347   0.10092787607256291   0.9493613198420622   0.5160845712704623   0.16188822575257056   0.742095120550388   0.16914459639432122   0.6221117905771991   0.036859750263745085   0.873763423095844   0.06139211381435736   0.812044503721134   0.19531677899718675   0.3293623977185131
0.6836340561003182   0.42493516871703746   0.19034848698367984   0.6785382296923688   0.9783291293187015   0.025349301612776255   0.31238172288100535   0.9830785949106174   0.6468141695664904   0.5252689166872071   0.10781790539297066   0.8821507188380545   0.6974528497244283   0.009184345416744885   0.9459296796404001   0.1400555982876665   0.5283082533301071   0.3870725548395458   0.909069929376655   0.2662921751918225   0.46691613951574973   0.5750280511184117   0.7137531503794683   0.9369297774733094   0.7832820834154315   0.1500928824013743   0.5234046633957884   0.2583915477809407   0.80495295409673   0.12474358078859804   0.21102294051478307   0.2753129528703233   0.15813878453023947   0.5994746641013909   0.10320503512181242   0.3931622340322688   0.46068593480581116   0.590290318684646   0.15727535548141233   0.2531066357446023   0.9323776814757041   0.20321776384510026   0.24820542610475732   0.9868144605527798   0.4654615419599543   0.6281897127266886   0.5344522757252891   0.04988468307947039   0.6821794585445229   0.4780968303253142   0.011047612329500611   0.7914931352985297   0.8772265044477929   0.35335324953671615   0.8000246718147175   0.5161801824282064   0.7190877199175535   0.7538785854353253   0.6968196366929051   0.12301794839593759   0.25840178511174233   0.16358826675067922   0.5395442812114928   0.8699113126513353
0.32602410363603823   0.9603705029055789   0.29133885510673546   0.8830968520985555   0.8605625616760839   0.33218079017889046   0.7568865793814464   0.8332121690190851   0.17838310313156105   0.8540839598535762   0.7458389670519457   0.04171903372055541   0.3011565986837681   0.50073071031686   0.9458142952372283   0.525538851292349   0.5820688787662146   0.7468521248815349   0.24899465854432315   0.4025209028964114   0.32366709365447227   0.5832638581308556   0.7094503773328303   0.5326095902450761   0.997642990018434   0.6228933552252767   0.41811152222609493   0.6495127381465207   0.1370804283423501   0.2907125650463862   0.6612249428446485   0.8163005691274355   0.9586973252107891   0.43662860519280994   0.9153859757927026   0.7745815354068801   0.657540726527021   0.9358978948759499   0.9695716805554744   0.24904268411453112   0.07547184776080636   0.1890457699944151   0.7205770220111513   0.8465217812181197   0.7518047541063341   0.6057819118635596   0.01112664467832091   0.31391219097304357   0.7541617640879   0.9828885566382829   0.593015122452226   0.6643994528265229   0.61708133574555   0.6921759915918967   0.9317901796075775   0.8480988836990874   0.6583840105347609   0.25554738639908675   0.016404203814874813   0.07351734829220723   0.0008432840077399598   0.3196494915231368   0.04683252325940038   0.8244746641776761
0.9253714362469336   0.1306037215287217   0.3262555012482491   0.9779528829595564   0.17356668214059953   0.5248218096651622   0.3151288565699282   0.6640406919865128   0.41940491805269947   0.5419332530268793   0.7221137341177022   0.9996412391599899   0.8023235823071495   0.8497572614349826   0.7903235545101247   0.15154235546090258   0.14393957177238859   0.594209875035896   0.7739193506952499   0.07802500716869536   0.14309628776464864   0.2745603835127591   0.7270868274358495   0.25355034299101925   0.21772485151771503   0.14395666198403737   0.40083132618760037   0.27559746003146285   0.044158169377115496   0.6191348523188751   0.0857024696176722   0.6115567680449501   0.6247532513244161   0.07720159929199581   0.36358873549997   0.61191552888496   0.8224296690172666   0.22744433785701318   0.5732651809898454   0.4603731734240575   0.678490097244878   0.6332344628211173   0.7993458302945955   0.38234816625536217   0.5353938094802293   0.3586740793083582   0.07225900285874597   0.1287978232643429   0.31766895796251426   0.21471741732432081   0.6714276766711456   0.8532003632328801   0.2735107885853988   0.5955825650054457   0.5857252070534734   0.24164359518793   0.6487575372609827   0.5183809657134498   0.22213647155350338   0.62972806630297   0.8263278682437163   0.2909366278564367   0.648871290563658   0.16935489287891242
0.14783777099883832   0.6577021650353194   0.8495254602690626   0.7870067266235503   0.612443961518609   0.2990280857269612   0.7772664574103166   0.6582089033592073   0.2947750035560947   0.08431066840264041   0.10583878073917104   0.8050085401263274   0.021264214970695933   0.48872810339719475   0.5201135736856977   0.5633649449383974   0.3725066777097132   0.9703471376837449   0.29797710213219425   0.9336368786354274   0.546178809465997   0.6794105098273082   0.6491058115685362   0.7642819857565151   0.3983410384671586   0.02170834479198878   0.7995803512994736   0.9772752591329648   0.7858970769485496   0.7226802590650275   0.022313893889157017   0.3190663557737574   0.4911220733924549   0.6383695906623872   0.916475113149986   0.51405781564743   0.469857858421759   0.1496414872651924   0.3963615394642883   0.9506928707090326   0.09735118071204578   0.17929434958144755   0.09838443733209407   0.017055992073605163   0.5511723712460489   0.49988383975413936   0.4492786257635578   0.2527740063170901   0.15283133277889024   0.47817549496215056   0.6496982744640842   0.2754987471841253   0.3669342558303406   0.755495235897123   0.6273843805749272   0.956432391410368   0.8758121824378857   0.11712564523473586   0.7109092674249412   0.44237457576293787   0.4059543240161268   0.9674841579695435   0.3145477279606529   0.49168170505390524
0.308603143304081   0.7881898083880959   0.21616329062855882   0.4746257129803001   0.7574307720580321   0.2883059686339566   0.766884664865001   0.22185170666320997   0.604599439279142   0.810130473671806   0.11718639040091676   0.9463529594790847   0.23766518344880128   0.054635237774683   0.4898020098259896   0.9899205680687168   0.36185300101091555   0.9375095925399471   0.7788927424010483   0.5475459923057789   0.9558986769947888   0.9700254345704037   0.4643450144403955   0.055864287251873646   0.6472955336907078   0.18183562618230778   0.24818172381183667   0.5812385742715735   0.8898647616326756   0.8935296575483512   0.4812970589468357   0.3593868676083636   0.2852653223535337   0.0833991838765452   0.36411066854591895   0.4130339081292789   0.04760013890473242   0.02876394610186219   0.8743086587199294   0.4231133400605621   0.6857471378938169   0.09125435356191505   0.09541591631888101   0.8755673477547833   0.7298484608990281   0.12122891899151135   0.6310709018784855   0.8197030605029096   0.08255292720832037   0.9393932928092036   0.38288917806664885   0.23846448623133604   0.19268816557564478   0.045863635260852374   0.9015921191198132   0.8790776186229725   0.9074228432221111   0.9624644513843071   0.5374814505738942   0.46604371049369353   0.8598227043173786   0.933700505282445   0.6631727918539648   0.042930370433131415
0.17407556642356176   0.84244615172053   0.5677568755350838   0.16736302267834816   0.44422710552453365   0.7212172327290186   0.9366859736565983   0.34765996217543854   0.3616741783162133   0.781823939919815   0.5537967955899494   0.10919547594410253   0.1689860127405685   0.7359603046589627   0.6522046764701364   0.23011785732113008   0.26156316951845743   0.7734958532746554   0.11472322589624212   0.7640741468274366   0.4017404652010788   0.8397953479922105   0.4515504340422773   0.7211437763943052   0.22766489877751703   0.9973491962716805   0.8837935585071934   0.5537807537159569   0.7834377932529833   0.27613196354266195   0.9471075848505952   0.20612079154051838   0.4217636149367701   0.4943080236228469   0.3933107892606457   0.09692531559641585   0.2527776021962016   0.7583477189638843   0.7411061127905094   0.8668074582752858   0.9912144326777442   0.9848518656892289   0.6263828868942672   0.10273331144784925   0.5894739674766654   0.14505651769701838   0.17483245285198995   0.38158953505354415   0.36180906869914836   0.14770732142533785   0.29103889434479646   0.8278087813375872   0.578371275446165   0.8715753578826759   0.3439313094942013   0.6216879897970689   0.15660766050939487   0.377267334259829   0.9506205202335556   0.524762674200653   0.9038300583131933   0.6189196152959446   0.20951440744304625   0.6579552159253672
0.9126156256354491   0.6340677496067159   0.583131520548779   0.555221904477518   0.32314165815878365   0.4890112319096975   0.40829906769678903   0.17363236942397384   0.9613325894596353   0.3413039104843596   0.11726017335199258   0.34582358808638664   0.3829613140134703   0.46972855260168367   0.7733288638577913   0.7241355982893177   0.2263536535040754   0.0924612183418547   0.8227083436242356   0.19937292408866478   0.3225235951908822   0.47354160304591003   0.6131939361811893   0.5414177081632976   0.4099079695554331   0.8394738534391941   0.030062415632410387   0.9861958036857795   0.08676631139664948   0.3504626215294967   0.6217633479356214   0.8125634342618058   0.12543372193701421   0.009158711045137095   0.5045031745836287   0.46673984617541914   0.742472407923544   0.5394301584434534   0.7311743107258375   0.7426042478861014   0.5161187544194685   0.4469689401015987   0.9084659671016019   0.5432313237974365   0.19359515922858633   0.9734273370556887   0.29527203092041243   0.0018136156341390169   0.7836871896731532   0.13395348361649453   0.2652096152880021   0.015617811948359445   0.6969208782765037   0.7834908620869978   0.6434462673523808   0.2030543776865537   0.5714871563394895   0.7743321510418607   0.138943092768752   0.7363145315111346   0.8290147484159456   0.23490199259840733   0.4077687820429145   0.9937102836250332
0.3128959939964771   0.7879330524968086   0.4993028149413127   0.45047895982759667   0.11930083476789077   0.8145057154411199   0.2040307840209002   0.44866534419345766   0.33561364509473757   0.6805522318246254   0.9388211687328981   0.43304753224509823   0.6386927668182338   0.8970613697376275   0.29537490138051736   0.22999315455854452   0.06720561047874432   0.1227292186957668   0.1564318086117654   0.49367862304740995   0.2381908620627987   0.8878272260973594   0.7486630265688509   0.4999683394223767   0.9252948680663217   0.09989417360055086   0.24936021162753824   0.04948937959478   0.8059940332984309   0.2853884581594309   0.04532942760663803   0.6008240354013223   0.47038038820369327   0.6048362263348056   0.1065082588737399   0.16777650315622414   0.8316876213854594   0.707774856597178   0.8111333574932225   0.9377833485976796   0.7644820109067151   0.5850456379014112   0.6547015488814572   0.4441047255502697   0.5262911488439164   0.6972184118040518   0.9060385223126063   0.944136386127893   0.6009962807775948   0.5973242382035009   0.656678310685068   0.894647006533113   0.7950022474791639   0.3119357800440699   0.6113488830784299   0.2938229711317907   0.32462185927547066   0.7070995537092644   0.5048406242046901   0.12604646797556654   0.49293423789001123   0.9993246971120864   0.6937072667114675   0.18826311937788692
0.7284522269832961   0.4142790592106751   0.03900571783001044   0.7441583938276172   0.20216107813937975   0.7170606474066233   0.1329671955174042   0.8000220076997242   0.601164797361785   0.11973640920312249   0.4762888848323362   0.9053750011666112   0.806162549882621   0.8078006291590526   0.8649400017539063   0.6115520300348205   0.4815406906071504   0.1007010754497882   0.36009937754921617   0.485505562059254   0.9886064527171392   0.10137637833770186   0.6663921108377486   0.29724244268136707   0.260154225733843   0.6870973191270268   0.6273863930077381   0.5530840488537498   0.05799314759446326   0.9700366717204033   0.494419197490334   0.7530620411540256   0.45682835023267826   0.8503002625172809   0.018130312657997767   0.8476870399874145   0.6506658003500572   0.0424996333582283   0.15319031090409155   0.23613500995259393   0.1691251097429068   0.9417985579084401   0.7930909333548753   0.75062944789334   0.18051865702576764   0.8404221795707383   0.12669882251712677   0.4533870052119729   0.9203644312919246   0.15332486044371152   0.4993124295093886   0.9003029563582231   0.8623712836974613   0.18328818872330818   0.004893232019054627   0.14724091520419744   0.4055429334647831   0.3329879262060273   0.9867629193610569   0.299553875216783   0.7548771331147259   0.29048829284779903   0.8335726084569653   0.06341886526418905
0.5857520233718191   0.3486897349393589   0.04048167510208995   0.3127894173708491   0.40523336634605145   0.5082675553686207   0.9137828525849632   0.8594024121588761   0.48486893505412687   0.3549426949249091   0.4144704230755746   0.9590994558006531   0.6224976513566655   0.17165450620160094   0.40957719105651996   0.8118585405964557   0.21695471789188242   0.8386665799955736   0.4228142716954631   0.5123046653796727   0.46207758477715655   0.5481782871477746   0.5892416632384978   0.4488858001154837   0.8763255614053375   0.19948855220841574   0.5487599881364078   0.13609638274463456   0.47109219505928596   0.6912209968397951   0.6349771355514446   0.27669397058575834   0.9862232600051591   0.33627830191488595   0.22050671247587006   0.31759451478510525   0.3637256086484936   0.164623795713285   0.8109295214193502   0.5057359741886496   0.1467708907566112   0.32595721571771136   0.388115249723887   0.9934313088089769   0.6846933059794547   0.7777789285699367   0.7988735864853892   0.5445455086934932   0.8083677445741172   0.578290376361521   0.2501135983489814   0.4084491259488586   0.33727554951483124   0.8870693795217259   0.6151364627975368   0.13175515536310026   0.35105228950967216   0.55079107760684   0.3946297503216667   0.814160640577995   0.9873266808611785   0.3861672818935549   0.5837002289023165   0.30842466638934546
0.8405557901045673   0.060210066175843575   0.19558497917842957   0.3149933575803686   0.1558624841251126   0.2824311376059068   0.39671139269304034   0.7704478488868755   0.34749473955099536   0.7041407612443858   0.14659779434405895   0.36199872293801677   0.010219190036164099   0.8170713817226599   0.5314613315465222   0.2302435675749165   0.659166900526492   0.26628030411582   0.13683158122485553   0.4160829269969215   0.6718402196653135   0.8801130222222651   0.553131352322539   0.10765826060757602   0.8312844295607462   0.8199029560464215   0.35754637314410936   0.7926649030272074   0.6754219454356336   0.5374718184405146   0.960834980451069   0.022217054140331965   0.3279272058846382   0.8333310571961288   0.81423718610701   0.6602183312023152   0.31770801584847413   0.01625967547346884   0.2827758545604878   0.42997476362739867   0.6585411153219821   0.7499793713576488   0.1459442733356323   0.013891836630477158   0.9867008956566686   0.8698663491353839   0.5928129210130934   0.9062335760229011   0.1554164660959225   0.049963393088962346   0.23526654786898404   0.11356867299569375   0.4799945206602889   0.5124915746484477   0.274431567417915   0.09135161885536178   0.15206731477565072   0.679160517452319   0.46019438131090495   0.4311332876530466   0.8343592989271766   0.6629008419788501   0.17741852675041714   0.001158524025647947
0.17581818360519447   0.9129214706212012   0.03147425341478481   0.9872666873951708   0.18911728794852578   0.04305512148581744   0.4386613324016914   0.08103311137226965   0.03370082185260328   0.9930917283968551   0.2033947845327074   0.9674644383765759   0.5537063011923143   0.48060015374840737   0.9289632171147924   0.8761128195212141   0.4016389864166636   0.8014396362960884   0.4687688358038874   0.4449795318681675   0.567279687489487   0.1385387943172383   0.29135030905347026   0.4438210078425196   0.39146150388429257   0.22561732369603704   0.25987605563868543   0.4565543204473488   0.20234421593576682   0.1825622022102196   0.821214723236994   0.37552120907507913   0.16864339408316353   0.18947047381336451   0.6178199387042866   0.4080567706985032   0.6149370928908492   0.7088703200649572   0.6888567215894943   0.5319439511772891   0.21329810647418554   0.9074306837688687   0.22008788578560687   0.08696441930912155   0.6460184189846985   0.7688918894516305   0.9287375767321366   0.6431434114666019   0.2545569151004059   0.5432745657555934   0.6688615210934512   0.18658909101925314   0.05221269916463911   0.3607123635453738   0.8476467978564572   0.811067881944174   0.8835693050814756   0.17124188973200927   0.22982685915217058   0.40301111124567074   0.2686322121906264   0.4623715696670521   0.5409701375626763   0.8710671600683817
0.055334105716440866   0.5549408858981834   0.32088225177706947   0.7841027407592601   0.40931568673174235   0.7860489964465529   0.39214467504493283   0.14095932929265817   0.15475877163133644   0.2427744306909595   0.7232831539514817   0.9543702382734051   0.10254607246669735   0.8820620671455857   0.8756363560950244   0.14330235632923102   0.21897676738522176   0.7108201774135764   0.6458094969428538   0.7402912450835603   0.9503445551945954   0.2484486077465243   0.10483935938017754   0.8692240850151786   0.8950104494781544   0.693507721848341   0.7839571076031081   0.08512134425591847   0.4856947627464121   0.9074587254017881   0.3918124325581752   0.9441620149632604   0.33093599111507566   0.6646842947108286   0.6685292786066936   0.9897917766898553   0.22838991864837832   0.7826222275652428   0.7928929225116692   0.8464894203606242   0.009413151263156547   0.07180205015166641   0.1470834255688153   0.10619817527706402   0.05906859606856118   0.8233534424051421   0.04224406618863775   0.23697409026188543   0.16405814659040668   0.12984572055680116   0.2582869585855297   0.15185274600596696   0.6783633838439945   0.22238699515501312   0.8664745260273544   0.20769073104270666   0.34742739272891887   0.5577027004441846   0.19794524742066083   0.21789895435285137   0.11903747408054058   0.7750804728789418   0.4050523249089917   0.3714095339922271
0.10962432281738403   0.7032784227272754   0.2579688993401764   0.26521135871516305   0.050555726748822846   0.8799249803221332   0.21572483315153865   0.02823726845327764   0.8864975801584162   0.7500792597653321   0.9574378745660089   0.8763845224473107   0.2081341963144216   0.5276922646103189   0.09096334853865455   0.668693791404604   0.8607068035855027   0.9699895641661345   0.8930181011179937   0.45079483705175266   0.7416693295049621   0.1949090912871927   0.48796577620900206   0.07938530305952558   0.6320450066875781   0.4916306685599174   0.22999687686882567   0.8141739443443625   0.5814892799387552   0.6117056882377842   0.01427204371728701   0.7859366758910848   0.6949916997803391   0.8616264284724521   0.056834169151278036   0.9095521534437742   0.4868575034659175   0.3339341638621331   0.9658708206126235   0.24085836203917016   0.6261506998804147   0.3639445996959987   0.07285271949462978   0.7900635249874175   0.8844813703754526   0.16903550840880596   0.5848869432856277   0.7106782219278919   0.25243636368787453   0.6774048398488887   0.3548900664168021   0.8965042775835294   0.6709470837491193   0.06569915161110448   0.3406180226995151   0.11056760169244452   0.9759553839687801   0.20407272313865243   0.28378385354823704   0.20101544824867032   0.4890978805028627   0.8701385592765194   0.3179130329356135   0.9601570862095001
0.8629471806224479   0.5061939595805207   0.24506031344098378   0.17009356122208266   0.9784658102469953   0.3371584511717147   0.660173370155356   0.45941533929419076   0.7260294465591207   0.6597536113228261   0.30528330373855395   0.5629110617106614   0.05508236281000149   0.5940544597117217   0.9646652810390389   0.45234346001821685   0.07912697884122132   0.3899817365730692   0.6808814274908018   0.2513280117695465   0.5900290983383586   0.5198431772965498   0.3629683945551883   0.29117092556004637   0.7270819177159107   0.01364921771602916   0.11790808111420456   0.12107736433796368   0.7486161074689154   0.6764907665443144   0.45773471095884855   0.6616620250437729   0.02258666090979466   0.016737155221488328   0.15245140722029457   0.09875096333311155   0.9675042980997932   0.42268269550976667   0.18778612618125565   0.6464075033148947   0.8883773192585719   0.03270095893669749   0.5069046986904537   0.39507949154534816   0.29834822092021324   0.5128577816401476   0.14393630413526545   0.10390856598530183   0.5712663032043025   0.4992085639241185   0.026028223021060885   0.9828312016473382   0.8226501957353871   0.822717797379804   0.5682935120622123   0.32116917660356525   0.8000635348255924   0.8059806421583157   0.4158421048419178   0.2224182132704537   0.8325592367257992   0.383297946648549   0.22805597866066216   0.576010709955559
0.9441819174672275   0.35059698771185155   0.7211512799702083   0.18093121841021081   0.6458336965470142   0.8377392060717039   0.577214975834943   0.07702265242490898   0.07456739334271167   0.33853064214758544   0.5511867528138821   0.09419145077757082   0.25191719760732456   0.5158128447677813   0.9828932407516696   0.7730222741740056   0.45185366278173217   0.7098322026094657   0.5670511359097519   0.5506040609035519   0.6192944260559329   0.3265342559609167   0.33899515724908974   0.9745933509479929   0.6751125085887055   0.9759372682490651   0.6178438772788813   0.7936621325377821   0.029278812041691298   0.13819806217736125   0.04062890144393844   0.7166394801128732   0.9547114186989796   0.7996674200297759   0.4894421486300564   0.6224480293353023   0.702794221091655   0.2838545752619945   0.5065489078783867   0.8494257551612967   0.2509405583099229   0.5740223726525288   0.9394977719686348   0.2988216942577448   0.63164613225399   0.24748811669161214   0.6005026147195451   0.32422834330975187   0.9565336236652845   0.271550848442547   0.9826587374406638   0.5305662107719697   0.9272548116235932   0.13335278626518576   0.9420298359967254   0.8139267306590967   0.9725433929246136   0.33368536623540995   0.45258768736666893   0.19147870132379438   0.26974917183295855   0.04983079097341548   0.9460387794882822   0.3420529461624977
0.01880861352303566   0.47580841832088666   0.006541007519647342   0.04323125190475289   0.3871624812690457   0.22832030162927452   0.4060383928001022   0.719002908595001   0.4306288576037612   0.9567694531867275   0.4233796553594384   0.1884366978230312   0.503374045980168   0.8234166669215417   0.48134981936271304   0.37450996716393453   0.5308306530555544   0.4897313006861318   0.028762131996044053   0.18303126584014015   0.2610814812225959   0.4399005097127163   0.08272335250776183   0.8409783196776425   0.24227286769956025   0.9640920913918296   0.07618234498811449   0.7977470677728896   0.8551103864305145   0.7357717897625551   0.6701439521880123   0.07874415917788857   0.4244815288267534   0.7790023365758276   0.24676429682857393   0.8903074613548574   0.9211074828465854   0.9555856696542858   0.7654144774658609   0.5157974941909228   0.3902768297910309   0.4658543689681541   0.7366523454698168   0.3327662283507827   0.129195348568435   0.02595385925543776   0.653928992962055   0.4917879086731402   0.8869224808688748   0.06186176786360812   0.5777466479739405   0.6940408409002506   0.03181209443836023   0.326089978101053   0.9076026957859282   0.6152966817223621   0.6073305656116069   0.5470876415252254   0.6608383989573543   0.7249892203675047   0.6862230827650215   0.5915019718709396   0.8954239214914934   0.2091917261765819
0.2959462529739906   0.12564760290278545   0.15877157602167652   0.8764254978257993   0.16675090440555557   0.0996937436473477   0.5048425830596215   0.384637589152659   0.2798284235366808   0.037831975783739584   0.927095935085681   0.6905967482524084   0.24801632909832055   0.7117419976826865   0.01949323929975272   0.07530006653004627   0.6406857634867137   0.16465435615746116   0.3586548403423984   0.35031084616254154   0.9544626807216922   0.5731523842865216   0.46323091885090506   0.14111911998595963   0.6585164277477016   0.44750478138373617   0.30445934282922854   0.2646936221601604   0.491765523342146   0.34781103773638844   0.799616759769607   0.8800560330075015   0.2119370998054652   0.30997906195264885   0.8725208246839261   0.18945928475509308   0.9639207707071447   0.5982370642699623   0.8530275853841733   0.1141592182250468   0.32323500722043097   0.4335827081125011   0.4943727450417749   0.7638483720625052   0.36877232649873876   0.8604303238259795   0.031141826190869897   0.6227292520765456   0.7102558987510372   0.41292554244224333   0.7266824833616413   0.3580356299163852   0.21849037540889119   0.06511450470585488   0.9270657235920343   0.47797959690888375   0.006553275603425982   0.755135442753206   0.05454489890810826   0.2885203121537907   0.04263250489628133   0.15689837848324373   0.2015173135239349   0.1743610939287439
0.7193974976758504   0.7233156703707426   0.70714456848216   0.41051272186623866   0.35062517117711156   0.8628853465447631   0.6760027422912901   0.787783469789693   0.6403692724260743   0.4499598041025198   0.9493202589296487   0.42974783987330784   0.4218788970171832   0.3848452993966649   0.022254535337614345   0.9517682429644241   0.41532562141375723   0.6297098566434589   0.9677096364295061   0.6632479308106334   0.3726931165174759   0.4728114781602152   0.7661923229055712   0.4888868368818895   0.6532956188416255   0.7494958077894726   0.059047754423411244   0.07837411501565084   0.3026704476645139   0.8866104612447094   0.38304501213212117   0.2905906452259578   0.6623011752384396   0.43665065714218965   0.4337247532024725   0.8608428053526499   0.24042227822125634   0.05180535774552474   0.41147021786485816   0.9090745623882258   0.8250966568074991   0.42209550110206584   0.4437605814353521   0.24582663157759246   0.4524035402900233   0.9492840229418507   0.6775682585297809   0.7569397946957029   0.7991079214483977   0.19978821515237816   0.6185205041063696   0.6785656796800521   0.4964374737838838   0.3131777539076687   0.23547549197424844   0.38797503445409437   0.8341362985454444   0.8765270967654791   0.8017507387717759   0.5271322291014444   0.593714020324188   0.8247217390199544   0.3902805209069178   0.6180576667132185
0.7686173635166889   0.4026262379178885   0.9465199394715657   0.37223103513562605   0.3162138232266656   0.45334221497603777   0.26895168094178484   0.6152912404399231   0.5171059017782678   0.2535539998236596   0.6504311768354152   0.9367255607598709   0.02066842799438397   0.9403762459159909   0.4149556848611668   0.5487505263057766   0.18653212944893968   0.0638491491505118   0.6132049460893909   0.021618297204332185   0.5928181091247517   0.23912741013055747   0.2229244251824731   0.4035606304911136   0.8242007456080629   0.836501172212669   0.27640448571090737   0.031329595355487586   0.5079869223813973   0.3831589572366312   0.007452804769122539   0.4160383549155645   0.9908810206031295   0.12960495741297157   0.35702162793370734   0.4793127941556936   0.9702125926087456   0.1892287114969807   0.9420659430725405   0.930562267849917   0.7836804631598059   0.12537956234646888   0.3288609969831497   0.9089439706455849   0.19086235403505417   0.8862521522159115   0.10593657180067657   0.5053833401544712   0.3666616084269913   0.04975098000324244   0.8295320860897692   0.4740537447989836   0.8586746860455939   0.6665920227666112   0.8220792813206467   0.05801538988341906   0.8677936654424644   0.5369870653536397   0.46505765338693933   0.5787025957277254   0.8975810728337189   0.347758353856659   0.5229917103143988   0.6481403278778085
0.11390060967391298   0.2223787915101901   0.19413071333124915   0.7391963572322237   0.9230382556388588   0.33612663929427866   0.08819414153057258   0.23381301707775248   0.5563766472118675   0.28637565929103626   0.2586620554408034   0.7597592722787689   0.6977019611662736   0.619783636524425   0.4365827741201567   0.7017438823953499   0.8299082957238092   0.08279657117078532   0.9715251207332174   0.12304128666762439   0.9323272228900903   0.7350382173141263   0.44853341041881856   0.4749009587898159   0.8184266132161773   0.5126594258039362   0.2544026970875694   0.7357046015575922   0.8953883575773185   0.17653278650965756   0.16620855555699685   0.5018915844798397   0.33901171036545097   0.8901571272186213   0.9075465001161934   0.7421323122010708   0.6413097491991774   0.27037349069419636   0.47096372599603675   0.04038842980572097   0.8114014534753682   0.18757691952341105   0.49943860526281936   0.9173471431380966   0.8790742305852779   0.4525387022092847   0.050905194844000794   0.4424461843482807   0.06064761736910062   0.9398792764053484   0.7965024977564313   0.7067415827906884   0.1652592597917821   0.7633464898956909   0.6302939421994346   0.20484999831084869   0.8262475494263312   0.8731893626770696   0.722747442083241   0.46271768610977787   0.18493780022715375   0.6028158719828732   0.25178371608720435   0.4223292563040569
0.37353634675178554   0.4152389524594622   0.752345110824385   0.5049821131659603   0.4944621161665076   0.9627002502501775   0.7014399159803842   0.06253592881767961   0.43381449879740697   0.022820973844829014   0.9049374182239528   0.35579434602699117   0.2685552390056249   0.25947448394913813   0.2746434760245183   0.15094434771614249   0.44230768957929373   0.38628512127206854   0.5518960339412772   0.6882266616063646   0.25736988935213995   0.7834692492891954   0.30011231785407283   0.26589740530230777   0.8838335426003544   0.3682302968297332   0.5477672070296878   0.7609152921363475   0.38937142643384687   0.4055300465795557   0.8463272910493036   0.6983793633186679   0.9555569276364398   0.38270907273472665   0.9413898728253508   0.3425850172916767   0.687001688630815   0.12323458878558856   0.6667463968008326   0.19164066957553422   0.24469399905152128   0.73694946751352   0.11485036285955538   0.5034140079691696   0.9873241096993813   0.9534802182243247   0.8147380450054825   0.23751660266686184   0.10349056709902688   0.5852499213945915   0.26697083797579474   0.47660131053051435   0.71411914066518   0.1797198748150358   0.4206435469264911   0.7782219472118465   0.7585622130287402   0.7970108020803092   0.4792536741011403   0.43563692992016984   0.07156052439792512   0.6737762132947206   0.8125072773003077   0.2439962603446356
0.8268665253464038   0.9368267457812005   0.6976569144407523   0.740582252375466   0.8395424156470225   0.9833465275568759   0.8829188694352698   0.5030656497086042   0.7360518485479957   0.3980966061622844   0.615948031459475   0.02646433917808983   0.021932707882815625   0.2183767313472486   0.19530448453298394   0.24824239196624331   0.2633704948540755   0.4213659292669395   0.7160508104318437   0.8126054620460735   0.19180997045615036   0.7475897159722189   0.903543533131536   0.5686092017014379   0.3649434451097465   0.8107629701910184   0.20588661869078367   0.8280269493259719   0.525401029462724   0.8274164426341425   0.3229677492555139   0.3249612996173677   0.7893491809147284   0.42931983647185806   0.7070197177960389   0.29849696043927787   0.7674164730319127   0.21094310512460945   0.511715233263055   0.05025456847303454   0.5040459781778373   0.78957717585767   0.7956644228312113   0.23764910642696102   0.3122360077216869   0.04198745988545106   0.8921208896996753   0.6690399047255231   0.9472925626119404   0.2312244896944327   0.6862342710088917   0.8410129553995512   0.42189153314921635   0.4038080470602902   0.3632665217533777   0.5160516557821835   0.632542352234488   0.9744882105884322   0.6562468039573388   0.21755469534290564   0.8651258792025752   0.7635451054638227   0.14453157069428382   0.1673001268698711
0.36107990102473797   0.9739679296061527   0.34886714786307255   0.92965102044291   0.048843893303051104   0.9319804697207017   0.4567462581633972   0.260611115717387   0.10155133069111073   0.700755980026269   0.7705119871545055   0.41959816031783576   0.6796597975418944   0.29694793296597877   0.4072454654011278   0.9035465045356522   0.04711744530740639   0.32245972237754655   0.750998661443789   0.6859918091927466   0.18199156610483114   0.5589146169137238   0.6064670907495051   0.5186916823228755   0.8209116650800932   0.584946687307571   0.2575999428864326   0.5890406618799654   0.772067771777042   0.6529662175868693   0.8008536847230354   0.32842954616257847   0.6705164410859313   0.9522102375606004   0.03034169756852989   0.9088313858447427   0.9908566435440369   0.6552623045946216   0.6230962321674021   0.00528488130909043   0.9437391982366305   0.3328025822170751   0.872097570723613   0.31929307211634383   0.7617476321317994   0.7738879653033512   0.26563047997410794   0.8006013897934683   0.9408359670517062   0.18894127799578014   0.008030537087675312   0.21156072791350292   0.1687681952746642   0.5359750604089107   0.2071768523646399   0.8831311817509244   0.4982517541887329   0.5837648228483103   0.17683515479610998   0.9742997959061818   0.507395110644696   0.9285025182536887   0.5537389226287079   0.9690149145970913
0.5636559124080655   0.5956999360366136   0.6816413519050948   0.6497218424807475   0.801908280276266   0.8218119707332624   0.4160108719309869   0.8491204526872792   0.8610723132245598   0.6328706927374823   0.4079803348433116   0.6375597247737763   0.6923041179498957   0.09689563232857151   0.2008034824786717   0.7544285430228518   0.19405236376116272   0.5131308094802611   0.023968327682561692   0.78012874711667   0.6866572531164667   0.5846282912265724   0.4702294050538538   0.8111138325195787   0.12300134070840132   0.9889283551899588   0.788588053148759   0.16139199003883117   0.3210930604321353   0.16711638445669647   0.3725771812177721   0.312271537351552   0.46002074720757546   0.5342456917192142   0.9645968463744605   0.6747118125777757   0.7677166292576799   0.4373500593906427   0.7637933638957889   0.9202832695549239   0.5736642654965172   0.9242192499103815   0.7398250362132271   0.1401545224382538   0.8870070123800504   0.339590958683809   0.26959563115937335   0.3290406899186751   0.7640056716716491   0.35066260349385014   0.4810075780106144   0.16764869987984393   0.44291261123951375   0.1835462190371537   0.1084303967928423   0.855377162528292   0.9828918640319383   0.6493005273179395   0.14383355041838178   0.18066534995051628   0.2151752347742584   0.21195046792729683   0.38004018652259297   0.2603820803955924
0.6415109692777412   0.2877312180169153   0.6402151503093658   0.12022755795733862   0.7545039568976909   0.9481402593331063   0.3706195191499924   0.7911868680386636   0.9904982852260418   0.5974776558392562   0.889611941139378   0.6235381681588196   0.547585673986528   0.4139314368021024   0.7811815443465358   0.7681610056305277   0.5646938099545897   0.7646309094841629   0.6373479939281539   0.5874956556800114   0.3495185751803313   0.5526804415568661   0.257307807405561   0.327113575284419   0.70800760590259   0.26494922353995076   0.6170926570961952   0.2068860173270803   0.9535036490048993   0.31680896420684446   0.24647313794620276   0.4156991492884168   0.9630053637788574   0.7193313083675883   0.3568611968068247   0.7921609811295972   0.4154196897923294   0.3053998715654859   0.575679652460289   0.023999975499069546   0.8507258798377397   0.540768962081323   0.9383316585321351   0.4365043198190582   0.5012073046574084   0.988088520524457   0.681023851126574   0.10939074453463922   0.7931996987548183   0.7231392969845062   0.06393119403037886   0.9025047272075589   0.8396960497499192   0.40633033277766173   0.8174580560841761   0.4868055779191421   0.8766906859710617   0.6869990244100734   0.4605968592773514   0.6946445967895449   0.4612709961787323   0.3815991528445875   0.8849172068170624   0.6706446212904753
0.6105451163409926   0.8408301907632645   0.9465855482849274   0.23414030147141718   0.10933781168358418   0.8527416702388075   0.2655616971583533   0.12474955693677796   0.3161381129287658   0.1296023732543014   0.20163050312797445   0.22224482972921908   0.47644206317884663   0.7232720404766397   0.3841724470437983   0.735439251810077   0.5997513772077849   0.0362730160665663   0.923575587766447   0.04079465502053206   0.13848038102905258   0.6546738632219788   0.03865838094938455   0.3701500337300567   0.52793526468806   0.8138436724587144   0.09207283266445719   0.13600973225863952   0.4185974530044758   0.9611020022199067   0.8265111355061039   0.01126017532186156   0.10245934007570999   0.8314996289656054   0.6248806323781294   0.7890153455926425   0.6260172768968634   0.10822758848896567   0.24070818533433108   0.053576093782565525   0.02626589968907845   0.07195457242239937   0.3171325975678841   0.012781438762033462   0.8877855186600259   0.41728070920042054   0.2784742166184996   0.6426314050319768   0.3598502539719659   0.6034370367417062   0.18640138395404238   0.5066216727733373   0.9412528009674901   0.6423350345217995   0.3598902484479385   0.4953614974514757   0.8387934608917801   0.8108354055561942   0.7350096160698091   0.7063461518588332   0.2127761839949168   0.7026078170672284   0.494301430735478   0.6527700580762676
0.18651028430583833   0.6306532446448291   0.17716883316759388   0.6399886193142342   0.29872476564581246   0.2133725354444085   0.8986946165490943   0.9973572142822574   0.9388745116738465   0.6099354987027023   0.712293232595052   0.4907355415089202   0.9976217107063564   0.9676004641809028   0.35240298414711346   0.9953740440574446   0.1588282498145763   0.1567650586247087   0.6173933680773044   0.28902789219861136   0.9460520658196595   0.4541572415574802   0.12309193734182637   0.6362578341223437   0.7595417815138212   0.8235039969126512   0.9459231041742324   0.9962692148081096   0.4608170158680087   0.6101314614682426   0.04722848762513814   0.998912000525852   0.5219425041941622   0.00019596276554035446   0.3349352550300862   0.5081764590169319   0.5243207934878058   0.03259549858463754   0.9825322708829727   0.5128024149594873   0.3654925436732294   0.8758304399599288   0.36513890280566835   0.223774522760876   0.4194404778535699   0.4216731984024486   0.242046965463842   0.5875166886385322   0.6598986963397487   0.5981692014897975   0.29612386128960955   0.5912474738304228   0.19908168047173996   0.9880377400215548   0.2488953736644714   0.5923354733045706   0.6771391762775778   0.9878417772560144   0.9139601186343852   0.08415901428763872   0.15281838278977203   0.9552462786713769   0.9314278477514124   0.5713565993281514
0.7873258391165426   0.07941583871144806   0.5662889449457441   0.34758207656727536   0.36788536126297267   0.6577426403089994   0.3242419794819021   0.7600653879287431   0.7079866649232239   0.05957343881920202   0.02811811819229257   0.16881791409832037   0.508904984451484   0.07153569879764722   0.7792227445278211   0.5764824407937498   0.8317658081739062   0.08369392154163278   0.8652626258934359   0.492323426506111   0.6789474253841342   0.1284476428702559   0.9338347781420235   0.9209668271779596   0.8916215862675916   0.04903180415880784   0.3675458331962794   0.5733847506106843   0.5237362250046189   0.3912891638498084   0.04330385371437734   0.8133193626819412   0.815749560081395   0.33171572503060637   0.015185735522084765   0.6445014485836208   0.30684457562991097   0.26018002623295916   0.23596299099426357   0.06801900778987106   0.4750787674560048   0.17648610469132636   0.3707003651008276   0.5756955812837601   0.7961313420718706   0.04803846182107047   0.43686558695880406   0.6547287541058004   0.9045097558042791   0.9990066576622626   0.06931975376252462   0.08134400349511611   0.3807735307996601   0.6077174938124542   0.02601590004814728   0.26802464081317495   0.5650239707182652   0.2760017687818479   0.010830164526062516   0.6235231922295541   0.25817939508835414   0.015821742548888722   0.7748671735317989   0.5555041844396831
0.7831006276323493   0.8393356378575624   0.40416680843097136   0.979808603155923   0.9869692855604787   0.7912971760364919   0.9673012214721673   0.32507984905012266   0.08245952975619973   0.7922905183742293   0.8979814677096427   0.24373584555500652   0.7016859989565396   0.184573024561775   0.8719655676614954   0.9757112047418316   0.13666202823827453   0.9085712557799271   0.8611354031354329   0.35218801251227744   0.8784826331499204   0.8927495132310383   0.08626822960363395   0.7966838280725944   0.09538200551757105   0.05341387537347604   0.6821014211726626   0.8168752249166713   0.1084127199570923   0.26211669933698417   0.7148001997004952   0.4917953758665487   0.025953190200892567   0.4698261809627549   0.8168187319908526   0.24805953031154218   0.32426719124435294   0.2852531564009799   0.9448531643293572   0.2723483255697106   0.1876051630060784   0.3766819006210528   0.08371776119392434   0.9201603130574332   0.309122529856158   0.4839323873900144   0.9974495315902904   0.12347648498483879   0.21374052433858695   0.43051851201653835   0.3153481104176278   0.30660126006816746   0.10532780438149467   0.16840181267955417   0.6005479107171325   0.8148058842016187   0.0793746141806021   0.6985756317167993   0.7837291787262799   0.5667463538900765   0.7551074229362492   0.41332247531581934   0.8388760143969226   0.29439802832036593
0.5675022599301708   0.03664057469476657   0.7551582532029983   0.37423771526293276   0.25837973007401277   0.5527081873047522   0.757708721612708   0.250761230278094   0.044639205735425805   0.12218967528821385   0.44236061119508013   0.9441599702099266   0.9393114013539311   0.9537878626086597   0.8418127004779477   0.1293540860083078   0.859936787173329   0.2552122308918604   0.058083521751667755   0.5626077321182312   0.10482936423707986   0.8418897555760411   0.2192075073547451   0.26820970379786535   0.5373271043069091   0.8052491808812745   0.46404925415174675   0.8939719885349325   0.27894737423289634   0.25254099357652227   0.7063405325390388   0.6432107582568386   0.23430816849747052   0.13035131828830843   0.2639799213439587   0.6990507880469121   0.2949967671435394   0.17656345567964873   0.42216722086601105   0.5696967020386042   0.43505997997021034   0.9213512247877883   0.3640836991143433   0.007088969920372974   0.33023061573313045   0.07946146921174731   0.1448761917595982   0.7388792661225076   0.7929035114262214   0.27421228833047284   0.6808269376078514   0.844907277587575   0.513956137193325   0.021671294753950576   0.9744864050688127   0.20169651933073643   0.2796479686958545   0.8913199764656422   0.7105064837248539   0.5026457312838244   0.9846512015523151   0.7147565207859934   0.28833926285884287   0.9329490292452202
0.5495912215821048   0.7934052959982051   0.9242555637444996   0.9258600593248472   0.21936060584897432   0.7139438267864577   0.7793793719849014   0.1869807932023395   0.4264570944227529   0.4397315384559849   0.09855243437704991   0.34207351561476446   0.9125009572294279   0.4180602437020343   0.12406602930823729   0.14037699628402805   0.6328529885335734   0.5267402672363922   0.41355954558338337   0.6377312650002037   0.6482017869812582   0.8119837464503987   0.12522028272454047   0.7047822357549836   0.0986105653991534   0.0185784504521937   0.2009647189800409   0.7789221764301364   0.879249959550179   0.30463462366573596   0.4215853469951395   0.5919413832277969   0.4527928651274261   0.864903085209751   0.3230329126180896   0.2498678676130324   0.5402919078979982   0.4468428415077167   0.19896688330985232   0.10949087132900436   0.9074389193644249   0.9201025742713245   0.785407337726469   0.4717596063288007   0.25923713238316665   0.10811882782092573   0.6601870550019285   0.7669773705738171   0.16062656698401326   0.08954037736873204   0.4592223360218876   0.9880551941436807   0.2813766074338342   0.7849057537029961   0.03763698902674807   0.3961138109158838   0.8285837423064081   0.9200026684932451   0.7146040764086584   0.14624594330285143   0.28829183440840983   0.4731598269855284   0.5156371930988062   0.036755071973847066
0.38085291504398494   0.5530572527142039   0.7302298553723372   0.5649954656450464   0.12161578266081831   0.4449384248932782   0.07004280037040872   0.7980180950712292   0.9609892156768051   0.3553980475245461   0.6108204643485211   0.8099629009275485   0.6796126082429709   0.5704922938215501   0.573183475321773   0.4138490900116647   0.8510288659365628   0.650489625328305   0.8585793989131146   0.2676031467088133   0.562737031528153   0.17732979834277657   0.3429422058143084   0.2308480747349662   0.18188411648416805   0.6242725456285727   0.6127123504419713   0.6658526090899198   0.060268333823349736   0.1793341207352945   0.5426695500715625   0.8678345140186906   0.09927911814654468   0.8239360732107484   0.9318490857230414   0.05787161309114203   0.4196665099035738   0.2534437793891983   0.3586656104012683   0.6440225230794773   0.568637643967011   0.6029541540608934   0.5000862114881537   0.376419376370664   0.005900612438857979   0.4256243557181168   0.15714400567384532   0.14557130163569781   0.82401649595469   0.8013518100895441   0.5444316552318741   0.479718692545778   0.7637481621313402   0.6220176893542496   0.0017621051603116   0.6118841785270874   0.6644690439847956   0.7980816161435013   0.06991301943727024   0.5540125654359453   0.24480253408122174   0.5446378367543029   0.7112474090360019   0.9099900423564681
0.6761648901142108   0.9416836826934095   0.2111611975478482   0.533570665985804   0.6702642776753528   0.5160593269752928   0.054017191874002904   0.38799936435010624   0.8462477817206628   0.7147075168857487   0.5095855366421288   0.9082806718043283   0.08249961958932263   0.09268982753149908   0.5078234314818172   0.2963964932772408   0.4180305756045271   0.29460821138799786   0.43791041204454695   0.7423839278412955   0.17322804152330537   0.749970374633695   0.726663003008545   0.8323938854848274   0.49706315140909463   0.8082866919402854   0.5155018054606968   0.29882321949902335   0.8267988737337418   0.2922273649649926   0.46148461358669396   0.9108238551489172   0.980551092013079   0.5775198480792438   0.9518990769445651   0.0025431833445889065   0.8980514724237564   0.4848300205477448   0.4440756454627479   0.7061466900673481   0.48002089681922927   0.19022180915974696   0.006165233418200935   0.9637627622260526   0.3067928552959239   0.44025143452605203   0.2795022304096559   0.13136887674122524   0.8097297038868293   0.6319647425857666   0.764000424948959   0.8325456572422019   0.9829308301530875   0.3397373776207741   0.30251581136226513   0.9217218020932848   0.0023797381400084655   0.7622175295415302   0.3506167344177   0.9191786187486959   0.10432826571625207   0.2773875089937854   0.9065410889549521   0.21303192868134777
0.6243073688970228   0.08716569983403846   0.9003758555367511   0.24926916645529512   0.3175145136010989   0.6469142653079865   0.6208736251270953   0.11790028971406988   0.5077848097142695   0.014949522722219756   0.8568732001781362   0.285354632471868   0.5248539795611821   0.6752121451014457   0.554357388815871   0.36363283037858324   0.5224742414211736   0.9129946155599155   0.20374065439817107   0.4444542116298874   0.4181459757049215   0.6356071065661301   0.29719956544321896   0.23142228294853964   0.7938386068078988   0.5484414067320915   0.3968237099064678   0.9821531164932445   0.47632409320679986   0.9015271414241052   0.7759500847793726   0.8642528267791746   0.9685392834925303   0.8865776187018853   0.9190768846012364   0.5788981943073066   0.44368530393134825   0.21136547360043972   0.3647194957853652   0.2152653639287234   0.9212110625101746   0.29837085804052427   0.16097884138719418   0.770811152298836   0.5030650868052531   0.6627637514743943   0.8637792759439752   0.5393888693502964   0.7092264799973543   0.1143223447423027   0.4669555660375074   0.5572357528570518   0.23290238679055447   0.21279520331819757   0.6910054812581349   0.6929829260778773   0.26436310329802415   0.3262175846163122   0.7719285966568985   0.1140847317705706   0.820677799366676   0.11485211101587245   0.4072091008715333   0.8988193678418472
0.8994667368565012   0.8164812529753481   0.2462302594843391   0.1280082155430112   0.39640165005124817   0.1537175015009539   0.3824509835403639   0.5886193461927148   0.6871751700538938   0.0393951567586512   0.9154954175028566   0.031383593335662964   0.45427278326333936   0.8265999534404537   0.22448993624472172   0.3384006672577857   0.18990967996531521   0.5003823688241414   0.4525613395878232   0.22431593548721512   0.3692318805986393   0.385530257808269   0.04535223871628995   0.32549656764536794   0.469765143742138   0.5690490048329209   0.7991219792319508   0.19748835210235674   0.0733634936908898   0.41533150333196694   0.41667099569158694   0.6088690059096419   0.38618832363699596   0.37593634657331576   0.5011755781887304   0.5774854125739789   0.9319155403736566   0.5493363931328621   0.2766856419440087   0.2390847453161932   0.7420058604083414   0.048954024308720666   0.8241243023561855   0.014768809828978073   0.3727739798097021   0.6634237665004517   0.7787720636398956   0.6892722421836102   0.9030088360675641   0.09437476166753081   0.9796500844079447   0.4917838900812534   0.8296453423766743   0.6790432583355639   0.5629790887163577   0.8829148841716115   0.44345701873967835   0.3031069117622481   0.06180351052762736   0.30542947159763256   0.5115414783660217   0.7537705186293859   0.7851178685836186   0.06634472628143935
0.7695356179576803   0.7048164943206653   0.9609935662274331   0.051575916452461276   0.3967616381479782   0.04139272782021364   0.1822215025875376   0.36230367426885113   0.4937528020804141   0.9470179661526829   0.20257141817959293   0.8705197841875978   0.6641074597037399   0.26797470781711896   0.6395923294632352   0.9876049000159862   0.22065044096406147   0.9648677960548709   0.5777888189356079   0.6821754284183537   0.7091089625980398   0.21109727742548495   0.7926709503519892   0.6158307021369144   0.9395733446403595   0.5062807831048196   0.8316773841245559   0.5642547856844531   0.5428117064923812   0.464888055284606   0.6494558815370184   0.2019511114156019   0.049058904411967114   0.5178700891319232   0.44688446335742543   0.33143132722800417   0.3849514447082273   0.2498953813148042   0.8072921338941903   0.34382642721201795   0.16430100374416584   0.2850275852599333   0.22950331495858245   0.6616509987936643   0.4551920411461261   0.07393030783444836   0.4368323646065933   0.045820296656749936   0.5156186965057666   0.5676495247296287   0.6051549804820373   0.4815655109722969   0.9728069900133854   0.10276146944502268   0.9556990989450189   0.279614399556695   0.9237480856014183   0.5848913803130995   0.5088146355875935   0.9481830723286908   0.538796640893191   0.3349959989982953   0.7015225016934032   0.6043566451166729
0.3744956371490252   0.049968413738361986   0.4720191867348208   0.9427056463230087   0.9193035960028991   0.9760381059039136   0.035186822128227505   0.8968853496662587   0.40368489949713243   0.4083885811742849   0.4300318416461902   0.41531983869396183   0.430877909483747   0.3056271117292622   0.4743327427011712   0.13570543913726682   0.5071298238823286   0.7207357314161628   0.9655181071135777   0.187522366808576   0.9683331829891376   0.38573973241786746   0.2639956054201744   0.5831657216919031   0.5938375458401124   0.3357713186795055   0.7919764186853536   0.6404600753688945   0.6745339498372133   0.35973321277559184   0.7567895965571261   0.7435747257026357   0.2708490503400809   0.9513446316013069   0.32675775491093595   0.32825488700867395   0.8399711408563338   0.6457175198720447   0.8524250122097647   0.19254944787140715   0.33284131697400526   0.924981788455882   0.8869069050961871   0.005027081062831154   0.36450813398486764   0.5392420560380145   0.6229112996760127   0.42186135937092806   0.7706705881447552   0.20347073735850904   0.830934880990659   0.7814012840020336   0.09613663830754193   0.8437375245829172   0.0741452844335329   0.0378265582993978   0.825287587967461   0.8923928929816103   0.747387529522597   0.7095716712907238   0.9853164471111272   0.24667537310956558   0.8949625173128323   0.5170222234193167
0.6524751301371219   0.32169358465368364   0.008055612216645244   0.5119951423564856   0.28796699615225424   0.7824515286156691   0.38514431254063264   0.09013378298555748   0.517296408007499   0.5789807912571601   0.5542094315499736   0.3087324989835239   0.42115976969995705   0.7352432666742429   0.48006414711644074   0.2709059406841261   0.595872181732496   0.8428503736926326   0.7326766175938437   0.5613342693934023   0.6105557346213688   0.596175000583067   0.8377141002810115   0.04431204597408558   0.9580806044842469   0.27448141592938347   0.8296584880643663   0.5323169036176001   0.6701136083319927   0.49202988731371433   0.4445141755237336   0.44218312063204257   0.1528172003244937   0.9130490960565543   0.8903047439737599   0.13345062164851867   0.7316574306245366   0.17780582938231132   0.41024059685731923   0.8625446809643925   0.1357852488920406   0.33495545568967866   0.6775639792634754   0.3012104115709903   0.5252295142706718   0.7387804551066116   0.839849878982464   0.2568983655969047   0.5671489097864248   0.46429903917722815   0.010191390918097771   0.7245814619793046   0.8970353014544321   0.9722691518635138   0.5656772153943642   0.2823983413472621   0.7442181011299385   0.059220055806959604   0.6753724714206042   0.14894771969874343   0.012560670505401814   0.8814142264246483   0.26513187456328496   0.28640303873435086
0.8767754216133612   0.5464587707349696   0.5875678952998095   0.9851926271633605   0.3515459073426895   0.807678315628358   0.7477180163173455   0.7282942615664558   0.7843969975562647   0.3433792764511298   0.7375266253992477   0.003712799587151195   0.8873616961018326   0.371110124587616   0.17184941000488352   0.721314458239889   0.1431435949718941   0.3118900687806564   0.4964769385842793   0.5723667385411456   0.13058292446649228   0.4304758423560081   0.23134506402099436   0.28596369980679476   0.2538075028531311   0.8840170716210385   0.6437771687211848   0.30077107264343417   0.9022615955104416   0.07633875599268052   0.8960591524038394   0.5724768110769783   0.11786459795417698   0.7329594795415507   0.15853252700459175   0.5687640114898271   0.23050290185234443   0.3618493549539347   0.9866831169997082   0.847449553249938   0.08735930688045034   0.04995928617327835   0.4902061784154289   0.27508281470879237   0.956776382413958   0.6194834438172703   0.25886111439443454   0.9891191149019977   0.702968879560827   0.7354663721962318   0.6150839456732496   0.6883480422585634   0.8007072840503854   0.6591276162035512   0.7190247932694102   0.1158712311815851   0.6828426860962084   0.9261681366620006   0.5604922662648185   0.547107219691758   0.45233978424386395   0.5643187817080658   0.5738091492651103   0.6996576664418199
0.3649804773634136   0.5143594955347874   0.08360297084968137   0.42457485173302756   0.40820409494945553   0.8948760517175173   0.8247418564552469   0.43545573683102995   0.7052352153886285   0.15940967952128546   0.2096579107819972   0.7471076945724665   0.9045279313382432   0.5002820633177342   0.490633117512587   0.6312364633908815   0.22168524524203484   0.5741139266557337   0.9301408512477686   0.08412924369912345   0.7693454609981709   0.009795144947667835   0.3563317019826583   0.3844715772573035   0.40436498363475726   0.4954356494128804   0.2727287311329769   0.959896725524276   0.9961608886853017   0.6005595976953632   0.4479868746777301   0.5244409886932461   0.2909256732966731   0.44114991817407767   0.23832896389573288   0.7773332941207796   0.3863977419584299   0.9408678548563434   0.7476958463831459   0.1460968307298981   0.1647124967163951   0.36675392820060976   0.8175549951353773   0.06196758703077466   0.39536703571822424   0.35695878325294195   0.46122329315271904   0.6774960097734711   0.9910020520834669   0.8615231338400616   0.18849456201974213   0.7175992842491952   0.9948411633981652   0.26096353614469847   0.740507687342012   0.19315829555594916   0.7039154901014921   0.8198136179706208   0.5021787234462792   0.41582500143516965   0.31751774814306216   0.8789457631142774   0.7544828770631333   0.26972817070527155
0.1528052514266671   0.5121918349136676   0.936927881927756   0.2077605836744969   0.7574382157084428   0.15523305166072565   0.4757045887750369   0.5302645739010258   0.7664361636249759   0.2937099178206641   0.2872100267552948   0.8126652896518306   0.7715950002268107   0.03274638167596563   0.5467023394132827   0.6195069940958814   0.06767951012531861   0.21293276370534484   0.04452361596700353   0.20368199266071174   0.7501617619822565   0.33398700059106745   0.2900407389038702   0.9339538219554402   0.5973565105555894   0.8217951656773999   0.3531128569761143   0.7261932382809433   0.8399182948471465   0.6665621140166742   0.8774082682010774   0.19592866437991754   0.07348213122217057   0.3728521961960101   0.5901982414457826   0.38326337472808697   0.30188713099535985   0.3401058145200445   0.0434959020324999   0.7637563806322055   0.23420762087004124   0.12717305081469968   0.9989722860654964   0.5600743879714938   0.4840458588877848   0.7931860502236322   0.7089315471616261   0.6261205660160536   0.8866893483321954   0.9713908845462323   0.3558186901855119   0.8999273277351103   0.04677105348504893   0.30482877052955815   0.4784104219844345   0.7039986633551928   0.9732889222628783   0.931976574333548   0.8882121805386519   0.3207352886271058   0.6714017912675185   0.5918707598135036   0.8447162785061519   0.5569789079949002
0.43719417039747727   0.46469770899880386   0.8457439924406556   0.9969045200234065   0.9531483115096925   0.6715116587751716   0.13681244527902947   0.3707839540073528   0.06645896317749704   0.7001207742289393   0.7809937550935176   0.47085662627224245   0.019687909692448116   0.39529200369938117   0.3025833331090831   0.7668579629170497   0.04639898742956975   0.46331542936583314   0.4143711525704312   0.4461226742899438   0.37499719616205124   0.8714446695523297   0.5696548740642793   0.8891437662950435   0.937803025764574   0.40674696055352577   0.7239108816236236   0.8922392462716371   0.9846547142548815   0.7352353017783542   0.5870984363445941   0.5214552922642843   0.9181957510773845   0.035114527549414846   0.8061046812510766   0.05059866599204188   0.8985078413849363   0.6398225238500337   0.5035213481419935   0.2837407030749923   0.8521088539553666   0.17650709448420052   0.08915019557156222   0.8376180287850484   0.4771116577933154   0.30506242493187086   0.519495321507283   0.948474262490005   0.5393086320287414   0.8983154643783451   0.7955844398836593   0.05623501621836784   0.5546539177738599   0.16308016259999092   0.2084860035390652   0.5347797239540836   0.6364581666964754   0.12796563505057607   0.4023813222879887   0.48418105796204164   0.737950325311539   0.4881431112005424   0.8988599741459953   0.2004403548870494
0.8858414713561724   0.3116360167163419   0.809709778574433   0.36282232610200094   0.4087298135628571   0.006573591784471029   0.29021445706715004   0.414348063611996   0.8694211815341157   0.10825812740612598   0.4946300171834907   0.35811304739362815   0.3147672637602558   0.945177964806135   0.2861440136444255   0.8233333234395446   0.6783090970637805   0.817212329755559   0.8837626913564368   0.339152265477503   0.9403587717522415   0.3290692185550166   0.9849027172104415   0.13871191059045357   0.054517300396069016   0.017433201838674722   0.17519293863600857   0.7758895844884527   0.645787486833212   0.010859610054203692   0.8849784815688585   0.36154152087645663   0.7763663052990962   0.9026014826480777   0.39034846438536785   0.0034284734828285016   0.4615990415388404   0.9574235178419427   0.1042044507409424   0.18009515004328389   0.78328994447506   0.14021118808638366   0.22044175938450558   0.8409428845657809   0.8429311727228185   0.8111419695313671   0.235539042174064   0.7022309739753274   0.7884138723267495   0.7937087676926924   0.06034610353805542   0.9263413894868747   0.14262638549353757   0.7828491576384886   0.17536762196919686   0.5647998686104181   0.3662600801944413   0.8802476749904109   0.785019157583829   0.5613713951275896   0.9046610386556009   0.9228241571484682   0.6808147068428866   0.3812762450843057
0.12137109418054094   0.7826129690620846   0.46037294745838103   0.5403333605185248   0.27843992145772245   0.9714709995307176   0.22483390528431701   0.8381023865431974   0.4900260491309729   0.1777622318380252   0.1644878017462616   0.9117609970563226   0.34739966363743535   0.3949130741995366   0.9891201797770647   0.3469611284459046   0.9811395834429941   0.5146653992091257   0.20410102219323573   0.785589733318315   0.07647854478739317   0.5918412420606574   0.5232863153503491   0.40431348823400937   0.9551074506068522   0.8092282729985728   0.06291336789196811   0.8639801277154846   0.6766675291491298   0.8377572734678552   0.8380794626076511   0.02587774117228717   0.18664148001815686   0.65999504162983   0.6735916608613894   0.11411674411596448   0.8392418163807215   0.2650819674302935   0.6844714810843248   0.7671556156700599   0.8581022329377275   0.7504165682211679   0.48037045889108904   0.9815658823517448   0.7816236881503342   0.15857532616051043   0.9570841435407399   0.5772523941177355   0.826516237543482   0.3493470531619376   0.8941707756487718   0.7132722664022509   0.14984870839435221   0.5115897796940824   0.05609131304112071   0.6873945252299638   0.9632072283761953   0.8515947380642522   0.38249965217973125   0.5732777811139993   0.12396541199547387   0.5865127706339588   0.6980281710954065   0.8061221654439394
0.2658631790577465   0.8360962024127909   0.21765771220431746   0.8245562830921945   0.4842394909074122   0.6775208762522805   0.26057356866357756   0.24730388897445904   0.6577232533639302   0.32817382309034293   0.36640279301480577   0.5340316225722082   0.507874544969578   0.8165840433962606   0.3103114799736851   0.8466370973422443   0.5446673165933826   0.9649893053320082   0.9278118277939539   0.2733593162282451   0.42070190459790874   0.3784765346980495   0.22978365669854736   0.4672371507843057   0.15483872554016226   0.5423803322852585   0.012125944494229893   0.6426808676921112   0.6705992346327501   0.864859456032978   0.7515523758306524   0.3953769787176521   0.01287598126881987   0.536685632942635   0.38514958281584655   0.861345356145444   0.5050014362992419   0.7201015895463745   0.0748381028421615   0.014708258803199658   0.9603341197058594   0.7551122842143663   0.14702627504820767   0.7413489425749545   0.5396322151079506   0.3766357495163168   0.9172426183496604   0.2741117917906489   0.38479348956778836   0.8342554172310582   0.9051166738554304   0.6314309240985377   0.7141942549350383   0.9693959611980802   0.15356429802477808   0.2360539453808856   0.7013182736662184   0.43271032825544514   0.7684147152089316   0.3747085892354416   0.1963168373669765   0.7126087387090706   0.69357661236677   0.36000033043224194
0.23598271766111717   0.9574964544947043   0.5465503373185624   0.6186513878572873   0.6963505025531666   0.5808607049783876   0.629307718968902   0.3445395960666385   0.31155701298537825   0.7466052877473293   0.7241910451134717   0.7131086719681008   0.59736275805034   0.777209326549249   0.5706267470886935   0.47705472658721515   0.8960444843841215   0.34449899829380387   0.802212031879762   0.10234613735177359   0.6997276470171451   0.6318902595847332   0.10863541951299195   0.7423458069195317   0.4637449293560279   0.6743938050900289   0.5620850821944295   0.1236944190622443   0.7673944268028613   0.09353310011164132   0.9327773632255275   0.7791548229956058   0.4558374138174831   0.34692781236431197   0.20858631811205594   0.06604615102750507   0.8584746557671431   0.5697184858150629   0.6379595710233624   0.5889914244402898   0.9624301713830216   0.22521948752125906   0.8357475391436004   0.4866452870885163   0.2627025243658765   0.5933292279365258   0.7271121196306085   0.7442994801689846   0.7989575950098485   0.9189354228464969   0.16502703743617894   0.6206050611067403   0.03156316820698726   0.8254023227348556   0.23224967421065137   0.8414502381111345   0.5757257543895041   0.4784745103705436   0.023663356098595427   0.7754040870836294   0.717251098622361   0.9087560245554807   0.385703785075233   0.18641266264333956
0.7548209272393395   0.6835365370342216   0.5499562459316325   0.6997673755548233   0.492118402873463   0.09020730909769578   0.822844126301024   0.9554678953858387   0.6931608078636144   0.17127188625119888   0.657817088864845   0.33486283427909824   0.6615976396566272   0.3458695635163433   0.4255674146541937   0.49341259616796374   0.08587188526712299   0.8673950531457997   0.4019040585555983   0.7180085090843343   0.36862078664476194   0.958639028590319   0.01620027348036529   0.5315958464409948   0.6137998594054225   0.27510249155609745   0.4662440275487328   0.8318284708861715   0.12168145653195943   0.18489518245840164   0.6433999012477087   0.8763605755003329   0.428520648668345   0.013623296207202769   0.9855828123828637   0.5414977412212346   0.7669230090117178   0.6677537326908595   0.56001539772867   0.04808514505327089   0.6810511237445949   0.8003586795450598   0.1581113391730717   0.3300766359689366   0.3124303370998329   0.8417196509547408   0.14191106569270642   0.7984807895279419   0.6986304776944104   0.5666171593986433   0.6756670381439737   0.9666523186417704   0.5769490211624511   0.3817219769402417   0.032267136896264884   0.09029174314143751   0.14842837249410604   0.3680986807330389   0.046684324513401196   0.5487940019202029   0.38150536348238817   0.7003449480421794   0.4866689267847312   0.500708856866932
0.7004542397377933   0.8999862684971196   0.3285575876116595   0.17063222089799537   0.3880239026379604   0.05826661754237885   0.1866465219189531   0.3721514313700535   0.6893934249435499   0.4916494581437355   0.5109794837749795   0.4054991127282831   0.11244440378109884   0.1099274812034938   0.47871234687871456   0.3152073695868456   0.9640160312869928   0.7418288004704549   0.43202802236531335   0.7664133676666427   0.5825106678046046   0.04148385242827541   0.9453590955805822   0.26570451079971075   0.8820564280668113   0.14149758393115577   0.6168015079689226   0.09507228990171536   0.4940325254288509   0.08323096638877692   0.43015498604996955   0.7229208585316619   0.804639100485301   0.5915815082450414   0.9191755022749901   0.31742174580337873   0.6921946967042022   0.48165402704154764   0.44046315539627556   0.0022143762165331583   0.7281786654172093   0.7398252265710927   0.008435133030962208   0.23580100854989045   0.14566799761260477   0.6983413741428174   0.06307603745038005   0.9700964977501797   0.2636115695457935   0.5568437902116616   0.4462745294814574   0.8750242078484644   0.7695790441169426   0.47361282382288467   0.01611954343148786   0.15210334931680247   0.9649399436316416   0.8820313155778432   0.09694404115649774   0.8346816035134237   0.27274524692743946   0.4003772885362956   0.6564808857602221   0.8324672272968906
0.5445665815102301   0.6605520619652029   0.64804575272926   0.5966662187470001   0.3988985838976253   0.9622106878223855   0.5849697152788799   0.6265697209968204   0.1352870143518318   0.4053668976107239   0.1386951857974225   0.751545513148356   0.3657079702348892   0.9317540737878393   0.12257564236593463   0.5994421638315536   0.40076802660324756   0.04972275820999601   0.025631601209436892   0.7647605603181299   0.12802277967580813   0.6493454696737004   0.36915071544921474   0.9322933330212393   0.583456198165578   0.9887934077084976   0.7211049627199547   0.3356271142742392   0.18455761426795278   0.026582719886112025   0.13613524744107486   0.7090573932774188   0.04927059991612097   0.6212158222753881   0.9974400616436524   0.9575118801290627   0.6835626296812318   0.6894617484875488   0.8748644192777177   0.3580697162975091   0.2827946030779842   0.6397389902775529   0.8492328180682809   0.5933091559793792   0.15477182340217605   0.9903935206038524   0.48008210261906614   0.6610158229581399   0.571315625236598   0.0016001128953549114   0.7589771398991114   0.32538870868390063   0.3867580109686452   0.9750173930092428   0.6228418924580366   0.6163313154064819   0.3374874110525242   0.35380157073385476   0.6254018308143842   0.6588194352774192   0.6539247813712925   0.6643398222463059   0.7505374115366664   0.3007497189799101
0.37113017829330824   0.024600831968753102   0.9013045934683855   0.7074405630005309   0.21635835489113223   0.034207311364900655   0.42122249084931945   0.04642474004239104   0.6450427296545342   0.032607198469545746   0.6622453509502081   0.7210360313584904   0.25828471868588904   0.05758980546030286   0.03940345849217156   0.1047047159520085   0.9207973076333649   0.7037882347264481   0.4140016276777874   0.4458852806745893   0.26687252626207236   0.03944841248014215   0.6634642161411209   0.14513556169467923   0.8957423479687641   0.014847580511389047   0.7621596226727354   0.43769499869414835   0.6793839930776319   0.9806402691464884   0.34093713182341595   0.3912702586517573   0.03434126342309763   0.9480330706769426   0.6786917808732079   0.6702342272932669   0.7760565447372085   0.8904432652166397   0.6392883223810363   0.5655295113412584   0.8552592371038438   0.1866550304901917   0.2252866947032489   0.11964423066666907   0.5883867108417714   0.14720661801004956   0.561822478562128   0.9745086689719898   0.6926443628730073   0.1323590374986605   0.7996628558893926   0.5368136702778415   0.013260369795375426   0.1517187683521721   0.45872572406597656   0.14554341162608422   0.9789191063722777   0.20368569767522948   0.7800339431927686   0.4753091843328173   0.20286256163506922   0.3132424324585897   0.1407456208117323   0.9097796729915589
0.34760332453122544   0.126587401968398   0.9154589261084833   0.7901354423248899   0.759216613689454   0.9793807839583485   0.3536364475463555   0.8156267733529   0.06657225081644676   0.847021746459688   0.5539735916569629   0.27881310307505847   0.053311881021071324   0.6953029781075158   0.09524786759098641   0.13326969144897424   0.07439277464879353   0.49161728043228636   0.31521392439821777   0.657960507116157   0.8715302130137244   0.17837484797369668   0.17446830358648546   0.748180834124598   0.5239268884824989   0.05178744600529868   0.25900937747800207   0.9580453917997082   0.7647102747930448   0.07240666204695023   0.9053729299316466   0.14241861844680823   0.6981380239765981   0.22538491558726229   0.35139933827468367   0.8636055153717498   0.6448261429555268   0.5300819374797464   0.25615147068369726   0.7303358239227755   0.5704333683067332   0.038464657047460084   0.9409375462854794   0.07237531680661856   0.6989031552930088   0.8600898090737634   0.766469242698994   0.3241944826820205   0.17497626681051   0.8083023630684647   0.507459865220992   0.3661490908823123   0.4102659920174652   0.7358957010215145   0.6020869352893453   0.2237304724355041   0.7121279680408672   0.5105107854342522   0.2506875970146617   0.36012495706375436   0.06730182508534044   0.9804288479545058   0.9945361263309644   0.6297891331409788
0.49686845677860725   0.9419641909070456   0.05359858004548499   0.5574138163343603   0.7979653014855984   0.08187438183328227   0.287129337346491   0.23321933365233977   0.6229890346750884   0.27357201876481757   0.779669472125499   0.8670702427700274   0.21272304265762312   0.537676317743303   0.17758253683615366   0.6433397703345234   0.5005950746167559   0.027165532309050836   0.926894939821492   0.28321481327076903   0.4332932495314155   0.046736684354545074   0.9323588134905275   0.6534256801297902   0.9364247927528082   0.10477249344749939   0.8787602334450425   0.09601186379542986   0.1384594912672099   0.022898111614217117   0.5916308960985515   0.8627925301430901   0.5154704565921215   0.7493260928493995   0.8119614239730525   0.9957222873730627   0.30274741393449844   0.21164977510609653   0.6343788871368988   0.3523825170385393   0.8021523393177425   0.18448424279704567   0.7074839473154069   0.06916770376777026   0.368859089786327   0.1377475584425006   0.7751251338248795   0.4157420236379801   0.4324342970335187   0.032975064995001226   0.896364900379837   0.3197301598425502   0.2939748057663088   0.010076953380784109   0.30473400428128544   0.4569376296994601   0.7785043491741872   0.2607508605313845   0.4927725803082329   0.4612153423263975   0.4757569352396888   0.049101085425288016   0.8583936931713341   0.10883282528785823
0.6736045959219463   0.8646168426282423   0.15090974585592717   0.03966512152008797   0.3047455061356193   0.7268692841857417   0.37578461203104774   0.6239230978821079   0.8723112091021006   0.6938942191907405   0.4794197116512108   0.30419293803955766   0.5783364033357917   0.6838172658099564   0.1746857073699254   0.8472553083400975   0.7998320541616045   0.42306640527857187   0.6819131270616925   0.3860399660137   0.3240751189219157   0.37396531985328385   0.8235194338903584   0.2772071407258418   0.6504705229999694   0.5093484772250415   0.6726096880344312   0.23754201920575382   0.3457250168643501   0.7824791930392998   0.2968250760033835   0.6136189213236459   0.4734138077622495   0.08858497384855929   0.8174053643521727   0.30942598328408827   0.8950774044264578   0.4047677080386029   0.6427196569822473   0.4621706749439908   0.09524535026485323   0.9817013027600311   0.9608065299205548   0.07613070893029075   0.7711702313429375   0.6077359829067472   0.13728709603019645   0.798923568204449   0.12069970834296816   0.09838750568170572   0.4646774079957652   0.5613815489986952   0.7749746914786181   0.31590831264240593   0.1678523319923817   0.9477626276750493   0.30156088371636863   0.22732333879384667   0.350446967640209   0.6383366443909609   0.4064834792899109   0.8225556307552437   0.7077273106579617   0.1761659694469702
0.31123812902505765   0.8408543279952126   0.7469207807374069   0.10003526051667942   0.5400678976821202   0.23311834508846546   0.6096336847072104   0.30111169231223045   0.419368189339152   0.13473083940675976   0.14495627671144518   0.7397301433135353   0.6443934978605339   0.8188225267643539   0.9771039447190635   0.7919675156384861   0.34283261414416527   0.5914991879705072   0.6266569770788545   0.1536308712475251   0.9363491348542544   0.7689435572152634   0.9189296664208928   0.9774649018005549   0.6251110058291968   0.9280892292200507   0.172008885683486   0.8774296412838756   0.08504310814707661   0.6949708841315853   0.5623752009762756   0.576317948971645   0.6656749188079246   0.5602400447248255   0.41741892426483046   0.8365878056581098   0.02128142094739078   0.7414175179604716   0.4403149795457669   0.044620290019623705   0.6784488068032255   0.14991832998996452   0.8136580024669124   0.8909894187720986   0.7420996719489712   0.3809747727747011   0.8947283360460196   0.9135245169715437   0.11698866611977442   0.45288554355465044   0.7227194503625336   0.03609487568766813   0.03194555797269781   0.7579146594230652   0.16034424938625802   0.45977692671602305   0.36627063916477315   0.19767461469823974   0.7429253251214276   0.6231891210579132   0.3449892182173824   0.4562570967377681   0.30261034557566063   0.5785688310382896
0.6665404114141569   0.3063387667478036   0.4889523431087482   0.687579412266191   0.9244407394651857   0.9253639939731024   0.5942240070627285   0.7740548952946473   0.8074520733454114   0.472478450418452   0.8715045567001949   0.7379600196069792   0.7755065153727135   0.7145637909953868   0.7111603073139369   0.27818309289095616   0.40923587620794033   0.516889176297147   0.9682349821925093   0.6549939718330429   0.06424665799055795   0.06063207955937898   0.6656246366168487   0.07642514079475327   0.3977062465764011   0.7542933128115754   0.17667229350810046   0.38884572852856225   0.47326550711121534   0.828929318838473   0.5824482864453719   0.6147908332339149   0.665813433765804   0.356450868420021   0.710943729745177   0.8768308136269357   0.8903069183930905   0.6418870774246342   0.9997834224312402   0.5986477207359795   0.48107104218515023   0.12499790112748714   0.03154844023873092   0.9436537489029366   0.4168243841945923   0.06436582156810816   0.3659238036218823   0.8672286081081834   0.019118137618191186   0.31007250875653275   0.18925151011378183   0.4783828795796211   0.5458526305069759   0.48114318991805977   0.6068032236684099   0.8635920463457062   0.8800391967411718   0.12469232149803876   0.8958594939232328   0.9867612327187705   0.9897322783480812   0.4828052440734046   0.8960760714919926   0.388113511982791
0.508661236162931   0.35780734294591743   0.8645276312532617   0.4444597630798543   0.09183685196833871   0.29344152137780927   0.49860382763137945   0.5772311549716709   0.07271871435014753   0.9833690126212765   0.3093523175175976   0.09884827539204978   0.5268660838431717   0.5022258227032168   0.7025490938491877   0.23525622904634355   0.646826887102   0.377533501205178   0.8066895999259549   0.24849499632757305   0.6570946087539187   0.8947282571317734   0.9106135284339621   0.860381484344782   0.14843337259098774   0.536920914185856   0.04608589718070044   0.4159217212649277   0.05659652062264902   0.24347939280804676   0.547482069549321   0.8386905662932568   0.9838778062725015   0.26011038018677024   0.23812975203172332   0.739842290901207   0.4570117224293298   0.7578845574835534   0.5355806581825356   0.5045860618548634   0.8101848353273299   0.38035105627837545   0.7288910582565807   0.25609106552729044   0.15309022657341115   0.48562279914660206   0.8182775298226185   0.3957095811825084   0.004656853982423416   0.948701884960746   0.772191632641918   0.9797878599175807   0.9480603333597744   0.7052224921526993   0.22470956309259713   0.14109729362432383   0.9641825270872729   0.44511211196592904   0.9865798110608738   0.40125500272311676   0.5071708046579431   0.6872275544823756   0.4509991528783382   0.8966689408682533
0.6969859693306132   0.3068764982040001   0.7221080946217575   0.6405778753409629   0.5438957427572021   0.8212536990573981   0.9038305647991389   0.24486829415845446   0.5392388887747787   0.8725518140966521   0.13163893215722083   0.2650804342408738   0.5911785554150043   0.16732932194395272   0.9069293690646237   0.12398314061654998   0.6269960283277314   0.7222172099780236   0.92034955800375   0.7227281378934333   0.11982522366978827   0.03498965549564809   0.46935040512541176   0.8260591970251799   0.422839254339175   0.728113157291648   0.7472423105036543   0.18548132168421708   0.8789435115819729   0.90685945823425   0.8434117457045154   0.9406130275257626   0.33970462280719427   0.03430764413759796   0.7117728135472945   0.6755325932848888   0.74852606739219   0.8669783221936452   0.8048434444826708   0.5515494526683388   0.12153003906445861   0.14476111221562157   0.8844938864789208   0.8288213147749056   0.001704815394670343   0.10977145671997349   0.4151434813535091   0.0027621177497256684   0.5788655610554954   0.38165829942832546   0.6679011708498548   0.8172807960655086   0.6999220494735223   0.4747988411940755   0.8244894251453394   0.876667768539746   0.3602174266663281   0.44049119705647755   0.11271661159804496   0.2011351752548572   0.6116913592741381   0.5735128748628323   0.30787316711537416   0.6495857225865184
0.49016132020967945   0.42875176264721077   0.42337928063645336   0.8207644078116128   0.48845650481500913   0.31898030592723725   0.008235799282944252   0.8180022900618872   0.9095909437595139   0.9373220064989117   0.3403346284330894   0.0007214939963785347   0.20966889428599148   0.4625231653048362   0.51584520328775   0.12405372545663254   0.8494514676196634   0.02203196824835867   0.40312859168970505   0.9229185502017754   0.23776010834552527   0.44851909338552637   0.09525542457433088   0.27333282761525696   0.7475987881358458   0.019767330738315603   0.6718761439378775   0.45256841980364415   0.25914228332083666   0.7007870248110784   0.6636403446549333   0.6345661297417571   0.34955133956132284   0.7634650183121666   0.32330571622184384   0.6338446357453785   0.1398824452753314   0.30094185300733034   0.8074605129340938   0.5097909102887459   0.290430977655668   0.27890988475897166   0.40433192124438877   0.5868723600869706   0.05267086931014272   0.8303907913734453   0.30907649667005793   0.3135395324717136   0.3050720811742969   0.8106234606351297   0.6372003527321803   0.8609711126680695   0.04592979785346024   0.10983643582405138   0.9735600080772471   0.22640498292631245   0.6963784582921374   0.34637141751188477   0.6502542918554033   0.592560347180934   0.556496013016806   0.045429564504554446   0.8427937789213094   0.08276943689218802
0.266065035361138   0.7665196797455828   0.43846185767692064   0.49589707680521744   0.2133941660509953   0.9361288883721375   0.1293853610068627   0.1823575443335038   0.9083220848766984   0.1255054277370077   0.49218500827468237   0.3213864316654343   0.8623922870232381   0.015668991912956315   0.5186250001974353   0.09498144873912186   0.16601382873110074   0.6692975744010715   0.868370708342032   0.5024211015581879   0.6095178157142948   0.623868009896517   0.025576929420722632   0.41965166466599985   0.34345278035315674   0.8573483301509343   0.5871150717438021   0.9237545878607825   0.13005861430216145   0.9212194417787969   0.4577297107369393   0.7413970435272786   0.22173652942546307   0.7957140140417892   0.965544702462257   0.42001061186184435   0.35934424240222496   0.7800450221288329   0.4469197022648217   0.3250291631227225   0.1933304136711242   0.11074744772776135   0.5785489939227897   0.8226080615645346   0.5838125979568295   0.48687943783124427   0.552972064502067   0.40295639689853474   0.24035981760367275   0.62953110768031   0.965856992758265   0.47920180903775234   0.1103012033015113   0.7083116659015131   0.5081272820213257   0.7378047655104737   0.8885646738760482   0.9125976518597239   0.5425825795590687   0.31779415364862934   0.5292204314738232   0.13255262973089102   0.09566287729424706   0.9927649905259068
0.33589001780269906   0.02180518200312968   0.5171138833714575   0.17015692896137222   0.7520774198458696   0.5349257441718854   0.9641418188693904   0.7672005320628374   0.5117176022421969   0.9053946364915755   0.9982848261111255   0.28799872302508517   0.40141639894068554   0.19708297059006236   0.4901575440897997   0.5501939575146115   0.5128517250646373   0.28448531873033844   0.947574964530731   0.2323998038659822   0.983631293590814   0.15193268899944745   0.8519120872364839   0.23963481334007536   0.6477412757881149   0.13012750699631775   0.3347982038650265   0.06947788437870313   0.8956638559422454   0.5952017628244324   0.3706563849956361   0.30227735231586567   0.3839462537000485   0.6898071263328569   0.3723715588845106   0.014278629290780463   0.9825298547593629   0.49272415574279455   0.8822140147947108   0.46408467177616897   0.4696781296947256   0.20823883701245607   0.9346390502639799   0.23168486791018675   0.48604683610391153   0.05630614801300863   0.08272696302749596   0.9920500545701114   0.8383055603157966   0.9261786410166909   0.7479287591624695   0.9225721701914082   0.9426417043735512   0.3309768781922585   0.3772723741668334   0.6202948178755426   0.5586954506735028   0.6411697518594016   0.004900815282322765   0.6060161885847621   0.5761655959141398   0.14844559611660704   0.12268680048761187   0.14193151680859323
0.10648746621941423   0.940206759104151   0.18804775022363196   0.9102466488984065   0.6204406301155027   0.8839006110911424   0.105320787196136   0.918196594328295   0.782135069799706   0.9577219700744515   0.35739202803366654   0.9956244241368868   0.8394933654261548   0.626745091882193   0.9801196538668331   0.37532960626134415   0.2807979147526521   0.9855753400227913   0.9752188385845104   0.769313417676582   0.7046323188385123   0.8371297439061843   0.8525320380968985   0.6273819008679887   0.598144852619098   0.8969229848020334   0.6644842878732665   0.7171352519695823   0.9777042225035953   0.013022373710891029   0.5591635006771305   0.7989386576412872   0.1955691527038893   0.05530040363643956   0.20177147264346398   0.8033142335044005   0.3560757872777345   0.4285553117542466   0.22165181877663087   0.4279846272430563   0.07527787252508239   0.4429799717314552   0.2464329801921205   0.6586712095664743   0.3706455536865701   0.6058502278252709   0.39390094209522203   0.031289308698485584   0.772500701067472   0.7089272430232375   0.7294166542219555   0.3141540567289033   0.7947964785638767   0.6959048693123465   0.17025315354482495   0.515215399087616   0.5992273258599874   0.6406044656759069   0.968481680901361   0.7119011655832156   0.24315153858225289   0.21204915392166035   0.7468298621247301   0.28391653834015934
0.1678736660571705   0.7690691821902051   0.5003968819326097   0.625245328773685   0.7972281123706004   0.16321895436493425   0.10649593983738762   0.5939560200751994   0.024727411303128326   0.4542917113416967   0.37707928561543214   0.2798019633462961   0.22993093273925166   0.7583868420293502   0.20682613207060715   0.76458656425868   0.6307036068792643   0.11778237635344327   0.23834445116924619   0.052685398675464415   0.38755206829701144   0.9057332224317829   0.49151458904451606   0.7687688603353051   0.21967840223984092   0.1366640402415778   0.9911177071119065   0.1435235315616201   0.42245028986924055   0.9734450858766436   0.8846217672745188   0.5495675114864207   0.3977228785661122   0.5191533745349468   0.5075424816590867   0.26976554814012454   0.16779194582686055   0.7607665325055967   0.30071634958847954   0.5051789838814446   0.5370883389475962   0.6429841561521533   0.06237189841923337   0.4524935852059801   0.14953627065058483   0.7372509337203704   0.5708573093747173   0.683724724870675   0.9298578684107439   0.6005868934787927   0.5797396022628108   0.5402011933090549   0.5074075785415034   0.6271418076021491   0.695117834988292   0.9906336818226342   0.10968469997539118   0.10798843306720221   0.18757535332920533   0.7208681336825097   0.9418927541485306   0.34722190056160557   0.8868590037407258   0.21568914980106513
0.40480441520093435   0.7042377444094522   0.8244871053214924   0.763195564595085   0.2552681445503495   0.9669868106890818   0.2536297959467751   0.07947083972441   0.3254102761396056   0.36639991721028914   0.6738901936839642   0.5392696464153551   0.8180026975981022   0.7392581096081401   0.9787723586956723   0.5486359645927209   0.7083179976227111   0.6312696765409379   0.7911970053664669   0.8277678309102112   0.7664252434741804   0.2840477759793323   0.9043380016257411   0.6120786811091461   0.36162082827324604   0.5798100315698801   0.07985089630424873   0.848883116514061   0.10635268372289651   0.6128232208807983   0.8262211003574736   0.7694122767896511   0.7809424075832909   0.2464233036705092   0.1523309066735094   0.23014263037429594   0.9629397099851886   0.5071651940623692   0.1735585479778372   0.681506665781575   0.2546217123624776   0.8758955175214312   0.38236154261137034   0.8537388348713639   0.48819646888829715   0.591847741542099   0.4780235409856292   0.2416601537622178   0.1265756406150511   0.012037709972218855   0.39817264468138047   0.39277703724815677   0.020222956892154614   0.39921448909142054   0.5719515443239068   0.6233647604585058   0.23928054930886372   0.15279118542091136   0.4196206376503974   0.3932221300842098   0.2763408393236751   0.6456259913585423   0.24606208967256024   0.7117154643026347
0.02171912696119748   0.769730473837111   0.8637005470611899   0.8579766294312708   0.5335226580729003   0.17788273229501206   0.3856770060755607   0.616316475669053   0.40694701745784917   0.16584502232279322   0.9875043613941802   0.22353943842089624   0.3867240605656946   0.7666305332313726   0.41555281707027336   0.6001746779623905   0.14744351125683083   0.6138393478104613   0.9959321794198759   0.20695254787818074   0.8711026719331557   0.9682133564519191   0.7498700897473157   0.495237083575546   0.8493835449719583   0.19848288261480806   0.8861695426861258   0.6372604541442752   0.315860886899058   0.020600150319796017   0.500492536610565   0.02094397847522221   0.9089138694412088   0.8547551279970028   0.5129881752163848   0.7974045400543259   0.5221898088755142   0.08812459476563014   0.09743535814611151   0.19722986209193547   0.3747462976186834   0.4742852469551688   0.1015031787262356   0.9902773142137548   0.5036436256855276   0.5060718905032497   0.3516330889789199   0.49504023063820873   0.6542600807135693   0.3075890078884417   0.4654635462927942   0.8577797764939336   0.33839919381451133   0.28698885756864567   0.9649710096822292   0.8368357980187113   0.42948532437330256   0.43223372957164286   0.45198283446584425   0.03943125796438532   0.9072955154977883   0.3441091348060127   0.3545474763197327   0.8422013958724498
0.5325492178791049   0.8698238878508439   0.2530442975934971   0.8519240816586952   0.028905592193577346   0.3637519973475941   0.9014112086145771   0.3568838510204864   0.374645511480008   0.05616298945915247   0.435947662321783   0.49910407452655287   0.03624631766549666   0.7691741318905068   0.4709766526395539   0.6622682765078416   0.6067609932921941   0.33694040231886396   0.018993818173709678   0.6228370185434563   0.6994654777944057   0.9928312675128512   0.664446341853977   0.7806356226710064   0.1669162599153008   0.12300737966200738   0.4114020442604798   0.9287115410123113   0.13801066772172343   0.7592553823144133   0.5099908356459026   0.5718276899918249   0.7633651562417154   0.7030923928552608   0.07404317332411964   0.07272361546527202   0.7271188385762187   0.9339182609647539   0.6030665206845657   0.4104553389574304   0.12035784528402467   0.59697785864589   0.5840727025108561   0.7876183204139742   0.42089236748961895   0.6041465911330387   0.9196263606568791   0.006982697742967729   0.25397610757431816   0.48113921147103134   0.5082243163963992   0.07827115673065642   0.11596543985259472   0.7218838291566181   0.9982334807504966   0.5064434667388314   0.3526002836108793   0.018791436301357323   0.924190307426377   0.4337198512735595   0.6254814450346605   0.08487317533660335   0.32112378674181125   0.023264512316129044
0.5051235997506359   0.48789531669071334   0.7370510842309552   0.23564619190215488   0.08423123226101693   0.8837487255576746   0.8174247235740761   0.22866349415918716   0.8302551246866988   0.4026095140866433   0.30920040717767683   0.15039233742853075   0.714289684834104   0.6807256849300252   0.3109669264271802   0.6439488706896992   0.3616894012232248   0.6619342486286679   0.3867766190008033   0.21022901941613978   0.7362079561885643   0.5770610732920645   0.06565283225899204   0.18696450710001072   0.23108435643792835   0.08916575660135113   0.3286017480280369   0.9513183151978558   0.14685312417691143   0.2054170310436765   0.5111770244539607   0.7226548210386686   0.3165979994902126   0.8028075169570332   0.2019766172762839   0.572262483610138   0.6023083146561086   0.12208183202700805   0.8910096908491036   0.9283136129204387   0.2406189134328838   0.4601475833983402   0.5042330718483004   0.7180845935042989   0.5044109572443196   0.8830865101062757   0.43858023958930836   0.5311200864042882   0.2733266008063912   0.7939207535049245   0.1099784915612715   0.5798017712064324   0.12647347662947978   0.588503722461248   0.5988014671073107   0.8571469501677637   0.8098754771392671   0.7856962055042148   0.39682484983102684   0.2848844665576257   0.2075671624831586   0.6636143734772068   0.5058151589819232   0.35657085363718705
0.9669482490502748   0.20346679007886656   0.001582087133622744   0.6384862601328881   0.4625372918059552   0.3203802799725909   0.5630018475443144   0.10736617372859997   0.18921069099956403   0.5264595264676663   0.4530233559830429   0.5275644025221676   0.06273721437008424   0.9379558040064182   0.8542218888757321   0.670417452354404   0.25286173723081706   0.1522595985022034   0.4573970390447053   0.3855329857967782   0.045294574747658495   0.48864522502499663   0.9515818800627822   0.028962132159591144   0.07834632569738369   0.2851784349461301   0.9499997929291595   0.390475872026703   0.6158090338914285   0.9647981549735393   0.38699794538484505   0.283109698298103   0.42659834289186443   0.4383386285058729   0.9339745894018021   0.7555452957759354   0.3638611285217802   0.5003828244994547   0.07975270052607002   0.08512784342153146   0.11099939129096312   0.34812322599725126   0.6223556614813647   0.6995948576247533   0.06570481654330462   0.8594780009722546   0.6707737814185826   0.6706327254651621   0.987358490845921   0.5742995660261245   0.7207739884894231   0.28015685343845914   0.3715494569544925   0.6095014110525853   0.33377604310457804   0.9970471551403561   0.944951114062628   0.17116278254671238   0.3998014537027759   0.24150185936442067   0.5810899855408478   0.6707799580472577   0.3200487531767059   0.15637401594288922
0.47009059424988475   0.32265673205000645   0.6976930916953412   0.456779158318136   0.40438577770658013   0.4631787310777518   0.026919310276758656   0.7861464328529738   0.41702728686065915   0.8888791650516273   0.30614532178733556   0.5059895794145147   0.045477829906166715   0.279377753999042   0.9723692786827575   0.5089424242741587   0.10052671584353869   0.10821497145232964   0.5725678249799816   0.26744056490973794   0.5194367303026909   0.43743501340507196   0.2525190718032757   0.11106654896684875   0.049346136052806126   0.1147782813550655   0.5548259801079345   0.6542873906487128   0.644960358346226   0.6515995502773136   0.5279066698311758   0.868140957795739   0.22793307148556685   0.7627203852256863   0.22176134804384032   0.3621513783812242   0.18245524157940013   0.48334263122664434   0.24939206936108282   0.8532089541070655   0.08192852573586144   0.37512765977431467   0.6768242443811012   0.5857683891973275   0.5624917954331706   0.9376926463692428   0.4243051725778255   0.47470184023047884   0.5131456593803645   0.8229143650141773   0.869479192469891   0.820414449581766   0.8681853010341385   0.1713148147368636   0.3415725226387151   0.9522734917860272   0.6402522295485716   0.40859442951117725   0.11981117459487482   0.5901221134048029   0.4577969879691715   0.925251798284533   0.8704191052337921   0.7369131592977374
0.37586846223331005   0.5501241385102182   0.1935948608526908   0.15114477010040975   0.8133766668001394   0.6124314921409755   0.7692896882748653   0.6764429298699309   0.300231007419775   0.7895171271267982   0.8998104958049743   0.8560284802881648   0.43204570638563655   0.6182023123899346   0.5582379731662591   0.9037549885021378   0.7917934768370649   0.2096078828787574   0.43842679857138434   0.31363287509733484   0.3339964888678934   0.28435608459422446   0.5680076933375923   0.5767197157995975   0.9581280266345834   0.7342319460840062   0.37441283248490154   0.4255749456991877   0.14475135983444393   0.12180045394303071   0.6051231442100362   0.7491320158292568   0.8445203524146689   0.33228332681623246   0.7053126484050619   0.8931035355410919   0.4124746460290324   0.7140810144262978   0.14707467523880283   0.9893485470389543   0.6206811691919675   0.5044731315475404   0.7086478766674185   0.6757156719416194   0.28668468032407407   0.22011704695331596   0.1406401833298262   0.09899595614202193   0.32855665368949066   0.48588510086930975   0.7662273508449247   0.6734210104428342   0.18380529385504674   0.364084646926279   0.16110420663488842   0.9242889946135774   0.3392849414403778   0.03180132011004656   0.4557915582298265   0.031185459072485475   0.9268102954113454   0.31772030568374876   0.3087168829910236   0.04183691203353125
0.30612912621937793   0.8132471741362083   0.6000690063236052   0.3661212400919118   0.019444445895303863   0.5931301271828924   0.45942882299377896   0.26712528394988994   0.6908877922058132   0.10724502631358263   0.6932014721488543   0.5937042735070557   0.5070824983507665   0.7431603793873036   0.5320972655139659   0.6694152788934783   0.16779755691038864   0.7113590592772571   0.0763057072841394   0.6382298198209928   0.24098726149904323   0.3936387535935083   0.7675888242931158   0.5963929077874616   0.9348581352796653   0.5803915794572999   0.1675198179695106   0.2302716676955497   0.9154136893843614   0.9872614522744075   0.7080909949757317   0.9631463837456598   0.22452589717854826   0.880016425960825   0.014889522826877338   0.36944211023860407   0.7174433988277819   0.13685604657352135   0.4827922573129115   0.7000268313451259   0.5496458419173932   0.4254969872962643   0.40648655002877204   0.06179701152413305   0.3086585804183499   0.03185823370275602   0.6388977257356563   0.4654041037366715   0.37380044513868466   0.45146665424545607   0.4713779077661457   0.23513243604112183   0.4583867557543232   0.4642052019710485   0.763286912790414   0.2719860522954621   0.2338608585757749   0.5841887760102236   0.7483973899635367   0.902543942056858   0.5164174597479931   0.44733272943670216   0.26560513265062524   0.20251711071173215
0.9667716178306   0.021835742140437868   0.8591185826218531   0.1407200991875991   0.6581130374122499   0.9899775084376818   0.2202208568861969   0.6753159954509276   0.2843125922735653   0.5385108541922258   0.7488429491200512   0.44018355940980575   0.8259258365192421   0.0743056522211773   0.9855560363296372   0.16819750711434367   0.5920649779434672   0.4901168762109538   0.23715864636610043   0.2656535650574857   0.07564751819547413   0.042784146774251595   0.9715535137154752   0.06313645434575357   0.10887590036487423   0.020948404633813728   0.112434931093622   0.9224163551581545   0.45076286295262424   0.030970896196131883   0.892214074207425   0.24710035970722694   0.16645027067905893   0.4924600420039061   0.1433711250873739   0.8069168002974212   0.34052443415981676   0.4181543897827288   0.15781508875773675   0.6387192931830775   0.7484594562163496   0.928037513571775   0.9206564423916364   0.3730657281255918   0.6728119380208755   0.8852533667975234   0.9491029286761611   0.3099292737798382   0.5639360376560012   0.8643049621637097   0.8366679975825392   0.38751291862168374   0.11317317470337693   0.8333340659675779   0.944453923375114   0.1404125589144568   0.946722904024318   0.3408740239636717   0.8010827982877401   0.3334957586170356   0.6061984698645012   0.9227196341809429   0.6432677095300033   0.6947764654339581
0.8577390136481516   0.9946821206091678   0.7226112671383671   0.3217107373083663   0.18492707562727623   0.10942875381164445   0.773508338462206   0.011781463528528088   0.6209910379712751   0.24512379164793474   0.9368403408796668   0.6242685449068444   0.5078178632678981   0.41178972568035693   0.9923864175045528   0.48385598599238755   0.5610949592435801   0.0709157017166852   0.1913036192168127   0.15036022737535193   0.9548964893790789   0.14819606753574227   0.5480359096868093   0.4555837619413938   0.09715747573092724   0.15351394692657439   0.8254246425484422   0.1338730246330275   0.912230400103651   0.04408519311492995   0.051916304086236244   0.1220915611044994   0.29123936213237595   0.7989614014669952   0.1150759632065694   0.49782301619765507   0.7834214988644779   0.3871716757866383   0.12268954570201661   0.013967030205267506   0.2223265396208977   0.3162559740699531   0.9313859264852039   0.8636068028299156   0.2674300502418188   0.16805990653421082   0.38335001679839464   0.4080230408885218   0.1702725745108916   0.014545959607636418   0.5579253742499525   0.2741500162554943   0.2580421744072406   0.9704607664927065   0.5060090701637162   0.1520584551509949   0.9668028122748646   0.17149936502571125   0.3909331069571468   0.6542354389533398   0.18338131341038677   0.7843276892390729   0.26824356125513016   0.6402684087480723
0.961054773789489   0.4680717151691199   0.33685763476992625   0.7766616059181568   0.6936247235476702   0.30001180863490906   0.9535076179715316   0.368638565029635   0.5233521490367786   0.2854658490272726   0.3955822437215792   0.09448854877414066   0.2653099746295381   0.31500508253456616   0.889573173557863   0.9424300936231458   0.29850716235467345   0.1435057175088549   0.4986400666007162   0.2881946546698059   0.1151258489442867   0.35917802826978196   0.230396505345586   0.6479262459217335   0.15407107515479765   0.891106313100662   0.8935388705756597   0.8712646400035768   0.46044635160712744   0.591094504465753   0.9400312526041281   0.5026260749739418   0.9370942025703488   0.30562865543848033   0.544449008882549   0.4081375261998012   0.6717842279408107   0.9906235729039141   0.654875835324686   0.4657074325766554   0.3732770655861372   0.8471178553950592   0.1562357687239698   0.17751277790684952   0.25815121664185053   0.48793982712527734   0.9258392633783837   0.529586531985116   0.1040801414870529   0.5968335140246153   0.03230039280272404   0.6583218919815391   0.6436337898799255   0.005739009558862244   0.09226914019859589   0.15569581700759724   0.7065395873095767   0.7001103541203819   0.5478201313160469   0.747558290807796   0.03475535936876598   0.7094867812164677   0.8929442959913609   0.28185085823114064
0.6614782937826288   0.8623689258214084   0.7367085272673911   0.10433808032429111   0.4033270771407782   0.37442909869613117   0.8108692638890074   0.5747515483391752   0.2992469356537253   0.7775955846715159   0.7785688710862834   0.9164296563576361   0.6556131457737998   0.7718565751126537   0.6862997308876874   0.7607338393500388   0.9490735584642231   0.07174622099227178   0.1384795995716405   0.01317554854224277   0.9143181990954572   0.36225943977580405   0.24553530358027956   0.7313246903111021   0.2528399053128284   0.4998905139543956   0.5088267763128884   0.626986609986811   0.8495128281720502   0.12546141525826443   0.697957512423881   0.05223506164763587   0.5502658925183249   0.3478658305867485   0.9193886413375978   0.1358054052899998   0.8946527467445251   0.5760092554740949   0.23308891044991034   0.375071565939961   0.9455791882803019   0.5042630344818231   0.09460931087826985   0.3618960173977182   0.031260989184844726   0.14200359470601903   0.8490740072979903   0.6305713270866161   0.7784210838720163   0.6421130807516234   0.3402472309851019   0.003584717099805022   0.928908255699966   0.5166516654933591   0.6422897185612209   0.9513496554521692   0.3786423631816412   0.16878583490661048   0.7229010772236231   0.8155442501621694   0.4839896164371161   0.5927765794325156   0.48981216677371275   0.44047268422220837
0.5384104281568142   0.08851354495069255   0.39520285589544285   0.07857666682449015   0.5071494389719695   0.9465099502446735   0.5461288485974526   0.4480053397378741   0.7287283550999532   0.30439686949305006   0.2058816176123507   0.4444206226380691   0.7998200993999871   0.7877452039996911   0.5635918990511298   0.49307096718589993   0.4211777362183459   0.6189593690930806   0.8406908218275068   0.6775267170237306   0.9371881197812298   0.02618278966056497   0.35087865505379406   0.23705403280152218   0.3987776916244156   0.9376692447098725   0.9556757991583512   0.15847736597703205   0.8916282526524462   0.9911592944651989   0.4095469505608986   0.710472026239158   0.16289989755249298   0.6867624249721488   0.2036653329485479   0.2660514036010889   0.3630797981525059   0.8990172209724577   0.6400734338974181   0.772980436415189   0.9419020619341599   0.28005785187937715   0.7993826120699112   0.09545371939145843   0.004713942152930107   0.2538750622188122   0.4485039570161172   0.8583996865899363   0.6059362505285145   0.3162058175089397   0.49282815785776607   0.6999223206129042   0.7143079978760684   0.3250465230437409   0.08328120729686744   0.9894502943737462   0.5514081003235753   0.638284098071592   0.8796158743483196   0.7233988907726573   0.18832830217106947   0.7392668770991343   0.23954244045090145   0.9504184543574683
0.2464262402369095   0.45920902521975715   0.44015982838099016   0.8549647349660099   0.2417122980839794   0.205333963000945   0.991655871364873   0.9965650483760736   0.6357760475554649   0.8891281454920053   0.49882771350710686   0.29664272776316947   0.9214680496793967   0.5640816224482644   0.4155465062102394   0.30719243338942326   0.37005994935582126   0.9257975243766724   0.5359306318619199   0.5837935426167659   0.18173164718475182   0.18653064727753804   0.29638819141101846   0.6333750882592976   0.9353054069478424   0.7273216220577808   0.8562283630300284   0.7784103532932877   0.6935931088638629   0.5219876590568359   0.8645724916651554   0.7818453049172139   0.05781706130839797   0.6328595135648306   0.3657447781580485   0.4852025771540445   0.13634901162900134   0.06877789111656625   0.950198271947809   0.17801014376462126   0.76628906227318   0.1429803667398939   0.4142676400858891   0.5942166011478554   0.5845574150884283   0.9564497194623558   0.11787944867487063   0.9608415128885578   0.6492520081405859   0.22912809740457496   0.2616510856448423   0.18243115959527012   0.955658899276723   0.7071404383477391   0.3970785939796869   0.40058585467805613   0.8978418379683251   0.07428092478290842   0.03133381582163844   0.9153832775240116   0.7614928263393237   0.005503033666342174   0.0811355438738294   0.7373731337593904
0.9952037640661436   0.8625226669264483   0.6668679037879403   0.14315653261153505   0.4106463489777154   0.9060729474640924   0.5489884551130696   0.18231501972297726   0.7613943408371294   0.6769448500595175   0.28733736946822735   0.9998838601277071   0.8057354415604064   0.9698044117117784   0.8902587754885404   0.599298005449651   0.9078936035920814   0.89552348692887   0.858924959666902   0.6839147279256393   0.14640077725275766   0.8900204532625279   0.7777894157930726   0.946541594166249   0.15119701318661402   0.027497786336079553   0.11092151200513227   0.8033850615547139   0.7405506642088986   0.1214248388719871   0.5619330568920626   0.6210700418317366   0.9791563233717692   0.4444799888124696   0.2745956874238353   0.6211861817040295   0.17342088181136275   0.4746755771006912   0.3843369119352949   0.02188817625437852   0.2655272782192814   0.5791520901718211   0.525411952268393   0.3379734483287392   0.11912650096652373   0.6891316369092934   0.7476225364753204   0.39143185416249027   0.9679294877799097   0.6616338505732138   0.6367010244701882   0.5880467926077764   0.22737882357101108   0.5402090117012267   0.0747679675781255   0.9669767507760397   0.2482225001992419   0.09572902288875706   0.8001722801542902   0.3457905690720103   0.07480161838787916   0.6210534457880659   0.4158353682189953   0.3239023928176318
0.8092743401685978   0.041901355616244716   0.8904234159506024   0.9859289444888926   0.690147839202074   0.3527697187069514   0.14280087947528192   0.5944970903264023   0.7222183514221643   0.6911358681337376   0.5060998550050938   0.006450297718625883   0.49483952785115326   0.15092685643251094   0.4313318874269683   0.039473546942586105   0.24661702765191135   0.055197833543753884   0.6311596072726781   0.6936829778705759   0.1718154092640322   0.434144387755688   0.2153242390536828   0.3697805850529441   0.36254106909543443   0.3922430321394433   0.3249008231030805   0.3838516405640515   0.6723932298933604   0.0394733134324919   0.18209994362779858   0.7893545502376492   0.9501748784711961   0.34833744529875427   0.6760000886227048   0.7829042525190233   0.45533535062004277   0.19741058886624335   0.24466820119573648   0.7434307055764372   0.20871832296813142   0.14221275532248945   0.6135085939230583   0.04974772770586141   0.03690291370409925   0.7080683675668015   0.39818435486937553   0.6799671426529174   0.6743618446086648   0.3158253354273582   0.07328353176629505   0.29611550208886583   0.001968614715304456   0.27635202199486625   0.8911835881384965   0.5067609518512166   0.05179373624410842   0.928014576696112   0.21518349951579172   0.7238566993321933   0.5964583856240656   0.7306039878298687   0.9705152983200552   0.980425993755756
0.3877400626559342   0.5883912325073791   0.3570067043969969   0.9306782660498947   0.350837148951835   0.8803228649405778   0.9588223495276214   0.25071112339697726   0.6764753043431702   0.5644975295132195   0.8855388177613263   0.9545956213081115   0.6745066896278656   0.28814550751835327   0.9943552296228297   0.4478346694568948   0.6227129533837572   0.3601309308222413   0.7791717301070381   0.7239779701247016   0.026254567759691618   0.6295269429923727   0.8086564317869828   0.7435519763689455   0.6385145051037574   0.04113571048499351   0.45164972738998593   0.8128737103190509   0.28767735615192247   0.1608128455444158   0.4928273778623646   0.5621625869220737   0.6112020518087523   0.5963153160311963   0.6072885601010383   0.6075669656139622   0.9366953621808867   0.308169808512843   0.6129333304782085   0.15973229615706735   0.3139824087971294   0.9480388776906017   0.8337616003711704   0.4357543260323658   0.28772784103743776   0.31851193469822897   0.025105168584187664   0.6922023496634203   0.6492133359336804   0.27737622421323543   0.5734554411942018   0.8793286393443693   0.3615359797817579   0.11656337866881965   0.08062806333183715   0.31716605242229573   0.7503339279730056   0.5202480626376234   0.4733395032307988   0.7095990868083336   0.8136385657921189   0.21207825412478046   0.8604061727525903   0.5498667906512662
0.49965615699498955   0.2640393764341788   0.026644572381419842   0.11411246461890046   0.2119283159575518   0.9455274417359498   0.0015394037972321763   0.4219101149554802   0.5627149800238714   0.6681512175227144   0.42808396260303044   0.5425814756111108   0.20117900024211352   0.5515878388538947   0.3474558992711933   0.22541542318881505   0.45084507226910797   0.03133977621627137   0.8741163960403945   0.5158163363804815   0.6372065064769891   0.819261522091491   0.013710223287804127   0.9659495457292152   0.13755034948199948   0.5552221456573121   0.9870656509063843   0.8518370811103148   0.9256220335244477   0.6096947039213623   0.9855262471091522   0.4299269661548346   0.3629070535005763   0.9415434863986478   0.5574422845061217   0.8873454905437238   0.16172805325846273   0.38995564754475304   0.2099863852349284   0.6619300673549087   0.7108829809893548   0.35861587132848166   0.335869989194534   0.14611373097442723   0.07367647451236575   0.5393543492369908   0.32215976590672984   0.180164185245212   0.9361261250303663   0.9841322035796787   0.3350941150003455   0.32832710413489724   0.010504091505918588   0.3744374996583164   0.34956786789119343   0.8984001379800626   0.6475970380053423   0.4328940132596686   0.7921255833850718   0.011054647436338863   0.48586898474687956   0.04293836571491555   0.5821391981501434   0.34912458008143016
0.7749860037575248   0.6843224943864339   0.24626920895560941   0.20301084910700293   0.701309529245159   0.1449681451494431   0.9241094430488795   0.022846663861790944   0.7651834042147928   0.16083594156976444   0.5890153280485341   0.6945195597268937   0.7546793127088741   0.786398441911448   0.2394474601573406   0.7961194217468311   0.10708227470353185   0.3535044286517794   0.44732187677226887   0.7850647743104923   0.6212132899566523   0.31056606293686384   0.8651826786221255   0.43594019422906205   0.8462272861991275   0.62624356855043   0.6189134696665161   0.23292934512205915   0.1449177569539684   0.4812754234009869   0.6948040266176365   0.2100826812602682   0.37973435273917566   0.32043948183122245   0.10578869856910246   0.5155631215333745   0.6250550400303014   0.5340410399197745   0.8663412384117618   0.7194436997865433   0.5179727653267696   0.18053661126799506   0.419019361639493   0.9343789254760512   0.8967594753701174   0.8699705483311312   0.5538366830173675   0.49843873124698906   0.05053218917098991   0.24372697978070124   0.9349232133508515   0.2655093861249299   0.9056144322170215   0.7624515563797143   0.24011918673321497   0.05542670486466172   0.5258800794778459   0.44201207454849184   0.1343304881641125   0.5398635833312873   0.9008250394475443   0.9079710346287174   0.26798924975235067   0.8204198835447438
0.3828522741207747   0.7274344233607223   0.8489698881128577   0.8860409580686928   0.48609279875065736   0.8574638750295911   0.2951332050954901   0.3876022268217037   0.43556060957966747   0.6137368952488899   0.36020999174463864   0.12209284069677376   0.5299461773626459   0.8512853388691756   0.1200908050114237   0.06666613583211205   0.0040660978848001145   0.4092732643206837   0.9857603168473112   0.5268025525008248   0.10324105843725574   0.5013022296919664   0.7177710670949605   0.7063826689560809   0.720388784316481   0.773867806331244   0.8688011789821029   0.8203417108873882   0.23429598556582362   0.9164039313016529   0.5736679738866127   0.4327394840656845   0.7987353759861562   0.302667036052763   0.21345798214197412   0.31064664336891074   0.2687891986235102   0.45138169718358745   0.09336717713055041   0.2439805075367987   0.2647231007387101   0.04210843286290375   0.10760686028323922   0.7171779550359739   0.16148204230145435   0.5408062031709374   0.38983579318827866   0.010795286079892972   0.44109325798497334   0.7669383968396934   0.5210346142061758   0.19045357519250478   0.20679727241914972   0.8505344655380406   0.947366640319563   0.7577140911268203   0.4080618964329935   0.5478674294852776   0.7339086581775889   0.4470674477579095   0.13927269780948331   0.0964857323016901   0.6405414810470385   0.20308694022111082
0.8745495970707732   0.054377299438786345   0.5329346207637993   0.4859089851851369   0.7130675547693188   0.5135710962678489   0.1430988275755206   0.4751136991052439   0.27197429678434554   0.7466326994281555   0.6220642133693448   0.28466012391273915   0.06517702436519582   0.8960982338901149   0.6746975730497818   0.5269460327859189   0.6571151279322023   0.34823080440483734   0.9407889148721928   0.07987858502800937   0.517842430122719   0.2517450721031473   0.3002474338251544   0.8767916448068985   0.6432928330519457   0.19736777266436092   0.7673128130613551   0.39088265962176166   0.9302252782826269   0.683796676396512   0.6242139854858345   0.9157689605165177   0.6582509814982813   0.9371639769683565   0.0021497721164897184   0.6311088366037785   0.5930739571330855   0.04106574307824164   0.3274521990667079   0.10416280381785964   0.9359588292008832   0.6928349386734043   0.38666328419451507   0.024284218789850265   0.4181163990781643   0.441089866570257   0.08641585036936066   0.1474925739829517   0.7748235660262185   0.2437220939058961   0.31910303730800554   0.7566099143611901   0.8445982877435917   0.5599254175093841   0.694889051822171   0.8408409538446724   0.1863473062453103   0.6227614405410276   0.6927392797056813   0.20973211724089383   0.5932733491122247   0.5816956974627859   0.36528708063897336   0.1055693134230342
0.6573145199113416   0.8888607587893816   0.9786237964444583   0.08128509463318394   0.23919812083317732   0.4477708922191246   0.8922079460750977   0.9337925206502322   0.4643745548069588   0.2040487983132285   0.5731049087670921   0.17718260628904217   0.6197762670633672   0.6441233808038445   0.8782158569449211   0.3363416524443698   0.4334289608180569   0.021361940262816875   0.18547657723923983   0.12660953520347595   0.8401556117058321   0.43966624280003097   0.8201894966002664   0.02104022178044175   0.1828410917944905   0.5508054840106493   0.8415657001558081   0.9397551271472578   0.9436429709613132   0.10303459179152474   0.9493577540807104   0.005962606497025587   0.4792684161543544   0.8989857934782962   0.37625284531361836   0.8287800002079835   0.8594921490909873   0.2548624126744518   0.4980369883686972   0.4924383477636136   0.4260631882729304   0.23350047241163494   0.31256041112945737   0.3658288125601377   0.5859075765670984   0.793834229611604   0.49237091452919096   0.3447885907796959   0.4030664847726078   0.2430287456009546   0.6508052143733828   0.40503346363243814   0.45942351381129465   0.13999415380942987   0.7014474602926724   0.3990708571354125   0.9801550976569402   0.24100836033113363   0.325194614979054   0.5702908569274291   0.12066294856595298   0.9861459476566818   0.8271576266103567   0.07785250916381548
0.6945997602930226   0.7526454752450469   0.5145972154808994   0.7120236966036778   0.10869218372592425   0.9588112456334429   0.02222630095170844   0.36723510582398183   0.7056256989533164   0.7157825000324883   0.3714210865783256   0.9622016421915437   0.24620218514202177   0.5757883462230584   0.6699736262856533   0.5631307850561311   0.26604708748508155   0.33477998589192476   0.34477901130659927   0.992839928128702   0.14538413891912857   0.34863403823524297   0.5176213846962425   0.9149874189648866   0.450784378626106   0.5959885629901961   0.0030241692153431376   0.2029637223612088   0.3420921949001817   0.6371773173567532   0.9807978682636347   0.835728616537227   0.6364664959468653   0.9213948173242649   0.6093767816853091   0.8735269743456833   0.39026431080484353   0.34560647110120646   0.9394031553996558   0.3103961892895521   0.12421722331976198   0.010826485209281698   0.5946241440930565   0.31755626116085   0.9788330844006334   0.6621924469740388   0.07700275939681396   0.4025688421959634   0.5280487057745274   0.06620388398384267   0.07397859018147082   0.19960511983475462   0.18595651087434567   0.4290265666270895   0.09318072191783612   0.36387650329752763   0.5494900149274804   0.5076317493028246   0.48380394023252704   0.4903495289518444   0.1592257041226368   0.16202527820161813   0.5444007848328712   0.17995333966229232
0.03500848080287484   0.15119879299233643   0.9497766407398148   0.8623970785014423   0.05617539640224142   0.4890063460182977   0.8727738813430008   0.45982823630547887   0.528126690627714   0.42280246203445504   0.79879529116153   0.26022311647072427   0.34217017975336833   0.9937758954073656   0.7056145692436939   0.8963466131731966   0.792680164825888   0.48614414610454093   0.22181062901116685   0.4059970842213522   0.6334544607032512   0.32411886790292277   0.6774098441782955   0.2260437445590599   0.5984459799003763   0.17292007491058636   0.7276332034384808   0.3636466660576176   0.5422705834981348   0.6839137288922886   0.8548593220954799   0.9038184297521387   0.014143892870420869   0.26111126685783365   0.056064030933949884   0.6435953132814144   0.6719737131170526   0.2673353714504681   0.350449461690256   0.7472487001082179   0.8792935482911646   0.7811912253459271   0.12863883267908913   0.3412516158868656   0.24583908758791345   0.45707235744300434   0.4512289885007935   0.11520787132780567   0.6473931076875371   0.28415228253241803   0.7235957850623128   0.7515612052701881   0.10512252418940228   0.6002385536401293   0.8687364629668328   0.8477427755180493   0.09097863131898141   0.33912728678229576   0.812672432032883   0.2041474622366349   0.41900491820192887   0.07179191533182766   0.462222970342627   0.4568987621284171
0.5397113699107643   0.2906006899859005   0.3335841376635379   0.11564714624155151   0.29387228232285084   0.8335283325428962   0.8823551491627444   0.00043927491374583846   0.6464791746353137   0.5493760500104782   0.15875936410043157   0.24887806964355777   0.5413566504459114   0.9491374963703487   0.29002290113359874   0.4011352941255084   0.45037801912693   0.6100102095880531   0.4773504691007157   0.1969878318888735   0.031373100925001104   0.5382182942562254   0.015127498758088732   0.7400890697604564   0.4916617310142368   0.24761760427032486   0.6815433610945508   0.6244419235189049   0.197789448691386   0.4140892717274287   0.7991882119318064   0.6240026486051591   0.5513102740560724   0.8647132217169506   0.6404288478313749   0.3751245789616013   0.009953623610160951   0.9155757253466018   0.3504059466977762   0.9739892848360928   0.559575604483231   0.3055655157585488   0.8730554775970605   0.7770014529472193   0.5282025035582298   0.7673472215023234   0.8579279788389718   0.03691238318676297   0.036540772543993044   0.5197296172319985   0.17638461774442088   0.41247045966785806   0.8387513238526071   0.10564034550456983   0.3771964058126144   0.788467811062699   0.2874410497965347   0.24092712378761924   0.7367675579812395   0.41334323210109775   0.27748742618637373   0.3253513984410174   0.3863616112834633   0.4393539472650049
0.7179118217031427   0.019785882682468614   0.5133061336864029   0.6623524943177855   0.1897093181449129   0.2524386611801452   0.6553781548474311   0.6254401111310225   0.15316854560091986   0.7327090439481466   0.4789935371030103   0.21296965146316446   0.3144172217483128   0.6270686984435768   0.10179713129039587   0.4245018404004654   0.02697617195177811   0.38614157465595755   0.3650295733091564   0.011158608299367668   0.7494887457654044   0.06079017621494014   0.9786679620256931   0.5718046610343628   0.03157692406226159   0.04100429353247153   0.46536182833929024   0.9094521667165772   0.8418676059173487   0.7885656323523264   0.8099836734918591   0.28401205558555476   0.6886990603164288   0.05585658840417971   0.33099013638884883   0.07104240412239028   0.37428183856811603   0.4287878899606029   0.22919300509845295   0.6465405637219249   0.34730566661633794   0.042646315304645355   0.8641634317892966   0.6353819554225572   0.5978169208509335   0.9818561390897053   0.8854954697636035   0.06357729438819441   0.566239996788672   0.9408518455572337   0.42013364142431325   0.15412512767161712   0.7243723908713233   0.15228621320490734   0.6101499679324541   0.8701130720860624   0.035673330554894425   0.09642962480072763   0.2791598315436053   0.7990706679636721   0.6613914919867784   0.6676417348401247   0.049966826445152365   0.15253010424174723
0.3140858253704405   0.6249954195354793   0.18580339465585582   0.51714814881919   0.716268904519507   0.6431392804457742   0.30030792489225233   0.45357085443099565   0.15002890773083497   0.7022874348885405   0.8801742834679391   0.29944572675937847   0.4256565168595117   0.5500012216836331   0.270024315535485   0.4293326546733161   0.38998318630461726   0.4535715968829055   0.9908644839918797   0.630261986709644   0.7285916943178389   0.7859298620427808   0.9408976575467273   0.4777318824678968   0.4145058689473984   0.16093444250730143   0.7550942628908714   0.9605837336487068   0.6982369644278914   0.5177951620615273   0.4547863379986192   0.5070128792177111   0.5482080566970565   0.8155077271729868   0.57461205453068   0.20756715245833257   0.12255153983754478   0.26550650548935373   0.30458773899519503   0.7782344977850165   0.7325683535329275   0.8119349086064482   0.3137232550033154   0.1479725110753725   0.003976659215088627   0.02600504656366741   0.37282559745658805   0.6702406286074757   0.5894707902676902   0.8650706040563659   0.6177313345657166   0.709656894958769   0.8912338258397988   0.3472754419948387   0.1629449965670974   0.20264401574105795   0.3430257691427423   0.5317677148218518   0.5883329420364174   0.9950768632827254   0.22047422930519753   0.26626120933249814   0.28374520304122236   0.2168423654977089
0.48790587577227   0.4543263007260499   0.970021948037907   0.06886985442233641   0.4839292165571814   0.42832125416238254   0.5971963505813189   0.39862922581486065   0.8944584262894911   0.5632506501060165   0.9794650160156023   0.6889723308560917   0.003224600449692373   0.21597520811117787   0.8165200194485049   0.48632831511503366   0.6601988313069501   0.6842074932893261   0.22818707741208755   0.4912514518323083   0.43972460200175256   0.4179462839568279   0.9444418743708652   0.2744090863345994   0.9518187262294825   0.963619983230778   0.9744199263329583   0.20553923191226298   0.46788950967230114   0.5352987290683955   0.3772235757516393   0.8069100060974023   0.57343108338281   0.972048078962379   0.3977585597360369   0.11793767524131069   0.5702064829331176   0.7560728708512011   0.581238540287532   0.631609360126277   0.9100076516261675   0.07186537756187503   0.3530514628754444   0.14035790829396871   0.470283049624415   0.6539190936050471   0.40860958850457924   0.8659488219593693   0.5184643233949324   0.690299110374269   0.43418966217162097   0.6604095900471063   0.05057481372263133   0.15500038130587357   0.056966086419981715   0.853499583949704   0.4771437303398214   0.1829523023434946   0.6592075266839448   0.7355619087083933   0.9069372474067038   0.4268794314922935   0.07796898639641284   0.1039525485821163
0.9969295957805363   0.3550140539304185   0.7249175235209684   0.9635946402881476   0.5266465461561213   0.7010949603253714   0.3163079350163892   0.09764581832877828   0.008182222761188813   0.010795849951102337   0.8821182728447682   0.43723622828167197   0.9576074090385575   0.8557954686452288   0.8251521864247865   0.5837366443319679   0.48046367869873613   0.6728431663017341   0.1659446597408417   0.8481747356235746   0.5735264312920323   0.24596373480944067   0.08797567334442886   0.7442221870414583   0.5765968355114961   0.8909496808790222   0.36305814982346046   0.7806275467533107   0.04995028935537482   0.18985472055365077   0.046750214807071235   0.6829817284245324   0.041768066594186005   0.17905887060254844   0.16463194196230302   0.24574550014286048   0.08416065755562853   0.3232634019573197   0.3394797555375165   0.6620088558108925   0.6036969788568924   0.6504202356555855   0.17353509579667484   0.8138341201873179   0.03017054756486007   0.4044565008461448   0.08555942245224597   0.0696119331458596   0.453573712053364   0.5135068199671227   0.7225012726287855   0.28898438639254886   0.4036234226979892   0.3236520994134719   0.6757510578217143   0.6060026579680164   0.36185535610380315   0.14459322881092346   0.5111191158594113   0.36025715782515594   0.27769469854817463   0.8213298268536038   0.17163936032189475   0.6982483020142634
0.6739977196912822   0.17090959119801835   0.9981042645252199   0.8844141818269455   0.6438271721264222   0.7664530903518736   0.9125448420729739   0.8148022486810859   0.19025346007305816   0.25294627038475087   0.19004356944418843   0.525817862288537   0.786630037375069   0.929294170971279   0.5142925116224741   0.9198152043205206   0.42477468127126583   0.7847009421603556   0.003173395763062859   0.5595580464953646   0.14707998272309122   0.9633711153067518   0.8315340354411681   0.8613097444811012   0.473082263031809   0.7924615241087334   0.8334297709159482   0.9768955626541557   0.8292550909053868   0.0260084337568599   0.9208849288429742   0.16209331397306984   0.6390016308323286   0.773062163372109   0.7308413593987858   0.6362754516845328   0.8523715934572597   0.84376799240083   0.21654884777631167   0.7164602473640124   0.4275969121859938   0.0590670502404744   0.2133754520132488   0.15690220086864773   0.28051692946290263   0.09569593493372264   0.3818414165720807   0.29559245638754655   0.8074346664310936   0.3032344108249892   0.5484116456561325   0.31869689373339083   0.9781795755257068   0.2772259770681293   0.6275267168131583   0.156603579760321   0.3391779446933781   0.5041638136960203   0.8966853574143725   0.5203281280757881   0.48680635123611843   0.6603958212951904   0.6801365096380608   0.8038678807117758
0.05920943905012461   0.6013287710547159   0.46676105762481196   0.6469656798431281   0.778692509587222   0.5056328361209933   0.08491964105273127   0.3513732234555816   0.9712578431561284   0.2023984252960041   0.5365079953965988   0.03267632972219072   0.9930782676304216   0.9251724482278748   0.9089812785834405   0.8760727499618697   0.6539003229370435   0.4210086345318545   0.012295921169067999   0.3557446218860816   0.16709397170092505   0.7606128132366642   0.3321594115310072   0.5518767411743057   0.10788453265080045   0.15928404218194825   0.8653983539061952   0.9049110613311776   0.3291920230635785   0.653651206060955   0.7804787128534639   0.5535378378755961   0.3579341799074501   0.45125278076495084   0.2439707174568652   0.5208615081534054   0.36485591227702846   0.5260803325370761   0.33498943887342475   0.6447887581915356   0.7109555893399849   0.10507169800522156   0.3226935177043567   0.28904413630545406   0.5438616176390599   0.3444588847685574   0.9905341061733495   0.7371673951311484   0.4359770849882595   0.18517484258660916   0.1251357522671543   0.8322563337999707   0.10678506192468103   0.5315236365256543   0.34465703941369036   0.27871849592437464   0.7488508820172309   0.08027085576070336   0.10068632195682514   0.7578569877709693   0.3839949697402025   0.5541905232236273   0.7656968830834004   0.11306822957943369
0.6730393804002175   0.44911882521840574   0.44300336537904367   0.8240240932739796   0.12917776276115756   0.10465994044984836   0.45246925920569414   0.08685669814283133   0.6932006777728981   0.9194850978632392   0.32733350693853985   0.2546003643428606   0.5864156158482171   0.38796146133758497   0.9826764675248495   0.975881868418486   0.8375647338309862   0.3076906055768816   0.8819901455680244   0.21802488064751668   0.45356976409078364   0.7535000823532543   0.11629326248462395   0.10495665106808298   0.7805303836905662   0.30438125713484854   0.6732898971055803   0.2809325577941033   0.6513526209294086   0.1997213166850002   0.2208206378998861   0.19407585965127203   0.9581519431565105   0.28023621882176103   0.8934871309613462   0.9394754953084113   0.3717363273082934   0.8922747574841761   0.9108106634364967   0.9635936268899254   0.5341715934773072   0.5845841519072944   0.028820517868472353   0.7455687462424088   0.08060182938652365   0.8310840695540401   0.9125272553838484   0.6406120951743257   0.30007144569595745   0.5267028124191915   0.23923735827826814   0.3596795373802224   0.6487188247665489   0.32698149573419133   0.018416720378382045   0.1656036777289504   0.6905668816100383   0.046745276912430314   0.1249295894170358   0.226128182420539   0.31883055430174495   0.1544705194282543   0.21411892598053908   0.2625345555306136
0.7846589608244376   0.5698863675209599   0.18529840811206674   0.5169658092882049   0.704057131437914   0.7388022979669198   0.27277115272821834   0.8763537141138791   0.40398568574195654   0.21209948554772828   0.033533794449950194   0.5166741767336567   0.7552668609754076   0.885117989813537   0.015117074071568148   0.3510704990047062   0.06469997936536927   0.8383727129011067   0.8901874846545323   0.12494231658416723   0.7458694250636243   0.6839021934728524   0.6760685586739933   0.8624077610535537   0.9612104642391867   0.11401582595189245   0.4907701505619265   0.34544195176534875   0.25715333280127267   0.37521352798497265   0.21799899783370819   0.4690882376514697   0.8531676470593161   0.16311404243724437   0.184465203383758   0.952414060917813   0.09790078608390852   0.27799605262370736   0.16934812931218984   0.6013435619131068   0.033200806718539255   0.4396233397226007   0.2791606446576575   0.47640124532893957   0.2873313816549149   0.7557211462497484   0.6030920859836643   0.6139934842753859   0.32612091741572824   0.6417053202978559   0.11232193542173774   0.26855153251003716   0.06896758461445554   0.2664917923128833   0.8943229375880296   0.7994632948585675   0.21579993755513938   0.1033777498756389   0.7098577342042716   0.8470492339407544   0.11789915147123085   0.8253816972519316   0.5405096048920818   0.24570567202764762
0.0846983447526916   0.3857583575293308   0.2613489602344242   0.769304426698708   0.7973669630977767   0.6300372112795825   0.65825687425076   0.1553109424233221   0.4712460456820484   0.9883318909817265   0.5459349388290222   0.886759409913285   0.4022784610675929   0.7218400986688432   0.6516120012409927   0.08729611505471746   0.18647852351245353   0.6184623487932044   0.9417542670367212   0.24024688111396303   0.06857937204122266   0.7930806515412728   0.4012446621446394   0.9945412090863154   0.9838810272885311   0.4073222940119421   0.13989570191021516   0.22523678238760736   0.1865140641907544   0.7772850827323596   0.4816388276594552   0.06992583996428527   0.7152680185087059   0.7889531917506332   0.935703888830433   0.18316643005100033   0.31298955744111306   0.06711309308178984   0.28409188758944026   0.09587031499628287   0.12651103392865953   0.4486507442885855   0.3423376205527191   0.8556234338823199   0.05793166188743687   0.6555700927473126   0.9410929584080797   0.8610822247960044   0.0740506345989058   0.24824779873537056   0.8011972564978646   0.635845442408397   0.8875365704081514   0.47096271600301093   0.3195584288384094   0.5659196024441118   0.17226855189944545   0.6820095242523778   0.3838545400079765   0.38275317239311146   0.8592789944583324   0.614896431170588   0.09976265241853623   0.28688285739682856
0.7327679605296729   0.1662456868820025   0.7574250318658171   0.43125942351450874   0.674836298642236   0.5106755941346899   0.8163320734577374   0.5701771987185044   0.6007856640433302   0.2624277953993193   0.015134816959872786   0.9343317563101072   0.7132490936351787   0.7914650793963084   0.6955763881214634   0.3684121538659955   0.5409805417357333   0.10945555514393057   0.3117218481134869   0.9856589814728841   0.681701547277401   0.49455912397334256   0.2119591956949507   0.6987761240760555   0.9489335867477281   0.3283134370913401   0.4545341638291336   0.26751670056154675   0.27409728810549205   0.8176378429566502   0.6382020903713962   0.6973395018430425   0.6733116240621618   0.5552100475573308   0.6230672734115235   0.7630077455329352   0.9600625304269831   0.7637449681610226   0.9274908852900601   0.3945955916669397   0.41908198869124974   0.654289413017092   0.6157690371765732   0.40893661019405564   0.7373804414138488   0.15973028904374934   0.40380984148162247   0.7101604861180001   0.7884468546661207   0.8314168519524092   0.9492756776524889   0.4426437855564534   0.5143495665606287   0.01377900899575905   0.31107358728109263   0.745304283713411   0.8410379424984669   0.4585689614384282   0.6880063138695691   0.9822965381804758   0.8809754120714838   0.6948239932774056   0.7605154285795092   0.5877009465135361
0.461893423380234   0.04053458026031373   0.14474639140293596   0.17876433631948044   0.7245129819663851   0.8808042912165643   0.7409365499213135   0.4686038502014803   0.9360661273002644   0.049387439264155134   0.7916608722688246   0.025960064645026936   0.42171656073963576   0.03560843026839609   0.48058728498773207   0.28065578093161603   0.580678618241169   0.5770394688299679   0.7925809711181628   0.29835924275114023   0.6997032061696852   0.8822154755525623   0.03206554253865376   0.7106582962376041   0.23780978278945125   0.8416808952922485   0.8873191511357178   0.5318939599181237   0.5132968008230661   0.9608766040756841   0.1463826012144043   0.06329010971664341   0.5772306735228016   0.911489164811529   0.35472172894557963   0.03733004507161647   0.15551411278316585   0.8758807345431329   0.8741344439578476   0.7566742641400005   0.5748354945419969   0.298841265713165   0.08155347283968471   0.4583150213888602   0.8751322883723116   0.41662579016060275   0.04948793030103095   0.747656725151256   0.6373225055828604   0.5749448948683542   0.16216877916531314   0.21576276523313234   0.12402570475979435   0.6140682907926701   0.015786177950908857   0.15247265551648895   0.5467950312369927   0.702579125981141   0.6610644490053292   0.11514261044487246   0.3912809184538269   0.8266983914380082   0.7869300050474817   0.358468346304872
0.8164454239118301   0.5278571257248432   0.705376532207797   0.9001533249160117   0.9413131355395183   0.11123133556424043   0.655888601906766   0.1524965997647557   0.303990629956658   0.5362864406958863   0.4937198227414528   0.9367338345316234   0.17996492519686366   0.9222181499032162   0.47793364479054395   0.7842611790151345   0.6331698939598709   0.21963902392207507   0.8168691957852148   0.669118568570262   0.241888975506044   0.3929406324840669   0.0299391907377331   0.31065022226538996   0.425443551594214   0.8650835067592237   0.32456265852993615   0.4104968973493782   0.4841304160546956   0.7538521711949833   0.6686740566231701   0.2580002975846225   0.18013978609803757   0.21756573049909705   0.17495423388171735   0.32126646305299916   0.00017486090117392388   0.2953475805958809   0.6970205890911734   0.5370052840378647   0.367004966941303   0.07570855667380585   0.8801513933059586   0.8678867154676028   0.125115991435259   0.682767924189739   0.8502122025682255   0.5572364932022128   0.699672439841045   0.8176844174305152   0.5256495440382893   0.14673959585283455   0.21554202378634946   0.06383224623553196   0.8569754874151192   0.8887392982682121   0.0354022376883119   0.846266515736435   0.6820212535334018   0.5674728352152129   0.03522737678713797   0.550918935140554   0.9850006644422284   0.030467551177348187
0.6682224098458349   0.47521037846674813   0.10484927113626984   0.16258083570974544   0.5431064184105759   0.7924424542770092   0.2546370685680443   0.6053443425075327   0.843433978569531   0.9747580368464939   0.728987524529755   0.45860474665469814   0.6278919547831814   0.9109257906109619   0.8720120371146358   0.5698654483864861   0.5924897170948695   0.06465927487452704   0.189990783581234   0.0023926131712731866   0.5572623403077316   0.513740339733973   0.20499011913900556   0.971925061993925   0.8890399304618967   0.0385299612672249   0.1001408480027357   0.8093442262841796   0.34593351205132067   0.24608750699021575   0.8455037794346913   0.20399988377664688   0.5024995334817898   0.27132947014372183   0.11651625490493642   0.7453951371219487   0.8746075786986083   0.36040367953275987   0.2445042177903006   0.17552968873546265   0.2821178616037388   0.2957444046582329   0.05451343420906662   0.17313707556418947   0.7248555212960072   0.7820040649242598   0.8495233150700611   0.20121201357026447   0.8358155908341106   0.7434741036570349   0.7493824670673254   0.3918677872860849   0.48988207878278994   0.49738659666681917   0.903878687632634   0.18786790350943805   0.9873825453010002   0.22605712652309734   0.7873624327276976   0.44247276638748934   0.11277496660239185   0.8656534469903374   0.5428582149373969   0.2669430776520267
0.8306571049986531   0.5699090423321046   0.4883447807283303   0.0938060020878372   0.10580158370264585   0.7879049774078448   0.6388214656582692   0.8925939885175728   0.26998599286853525   0.04443087375080987   0.8894389985909439   0.5007262012314878   0.7801039140857453   0.5470442770839907   0.9855603109583099   0.31285829772204976   0.7927213687847452   0.32098715056089333   0.19819787823061236   0.8703855313345604   0.6799464021823532   0.4553337035705559   0.6553396632932155   0.6034424536825338   0.8492892971837003   0.8854246612384513   0.1669948825648851   0.5096364515946966   0.7434877134810544   0.09751968383060651   0.5281734169066158   0.6170424630771238   0.4735017206125191   0.05308881007979664   0.6387344183156719   0.11631626184563607   0.6933978065267739   0.506044532995806   0.653174107357362   0.8034579641235863   0.9006764377420287   0.1850573824349126   0.4549762291267497   0.9330724327890259   0.22073003555967535   0.7297236788643567   0.7996365658335343   0.32962997910649205   0.37144073837597513   0.8442990176259054   0.6326416832686491   0.8199935275117954   0.6279530248949208   0.7467793337952989   0.10446826636203334   0.20295106443467156   0.1544513042824016   0.6936905237155022   0.4657338480463614   0.0866348025890355   0.4610534977556278   0.18764599071969632   0.8125597406889994   0.2831768384654492
0.5603770600135992   0.0025886082847837106   0.3575835115622497   0.35010440567642337   0.3396470244539238   0.272864929420427   0.5579469457287155   0.02047442656993134   0.9682062860779487   0.42856591179452164   0.9253052624600663   0.2004808990581359   0.34025326118302796   0.6817865779992227   0.820836996098033   0.9975298346234643   0.18580195690062634   0.9880960542837205   0.3551031480516716   0.9108950320344289   0.7247484591449985   0.8004500635640242   0.5425434073626721   0.6277181935689796   0.16437139913139936   0.7978614552792405   0.1849598958004225   0.27761378789255625   0.8247243746774755   0.5249965258588134   0.627012950071707   0.25713936132262494   0.8565180885995268   0.09643061406429183   0.7017076876116407   0.056658462264489035   0.5162648274164989   0.4146440360650691   0.8808706915136078   0.05912862764102468   0.3304628705158726   0.4265479817813486   0.5257675434619361   0.14823359560659582   0.605714411370874   0.6260979182173244   0.983224136099264   0.5205154020376161   0.4413430122394747   0.828236462938084   0.7982642402988415   0.2429016141450599   0.6166186375619992   0.30323993707927055   0.17125129022713445   0.985762252822435   0.7601005489624723   0.2068093230149787   0.46954360261549377   0.9291037905579459   0.24383572154597338   0.7921652869499096   0.588672911101886   0.8699751629169212
0.9133728510301008   0.36561730516856095   0.06290536763994994   0.7217415673103255   0.30765843965922673   0.7395193869512365   0.07968123154068603   0.20122616527270923   0.8663154274197521   0.9112829240131525   0.2814169912418446   0.9583245511276494   0.2496967898577529   0.6080429869338819   0.11016570101471014   0.9725622983052143   0.4895962408952806   0.40123366391890325   0.6406220983992164   0.04345850774726844   0.24576051934930723   0.6090683769689936   0.05194918729733033   0.1734833448303472   0.3323876683192064   0.24345107180043268   0.9890438196573804   0.45174177752002176   0.024729228659979664   0.5039316848491961   0.9093625881166943   0.25051561224731256   0.1584138012402276   0.5926487608360437   0.6279455968748497   0.2921910611196632   0.9087170113824747   0.9846057739021616   0.5177798958601396   0.31962876281444885   0.4191207704871941   0.5833721099832584   0.8771577974609233   0.2761702550671804   0.1733602511378869   0.9743037330142648   0.8252086101635929   0.1026869102368332   0.8409725828186805   0.7308526612138321   0.8361647905062125   0.6509451327168114   0.8162433541587009   0.2269209763646359   0.9268022023895182   0.40042952046949887   0.6578295529184732   0.6342722155285923   0.2988566055146684   0.10823845934983568   0.7491125415359985   0.6496664416264305   0.7810767096545288   0.7886096965353868
0.32999177104880434   0.06629433164317212   0.9039189121936055   0.5124394414682064   0.15663151991091748   0.09199059862890734   0.07871030203001257   0.40975253123137323   0.31565893709223697   0.36113793741507527   0.24254551152380002   0.7588073985145618   0.49941558293353616   0.13421696105043934   0.31574330913428184   0.35837787804506294   0.8415860300150629   0.4999447455218471   0.016886703619613468   0.25013941869522727   0.0924734884790645   0.8502783038954166   0.2358099939650847   0.46152972215984045   0.7624817174302602   0.7839839722522444   0.33189108177147925   0.9490902806916339   0.6058501975193427   0.6919933736233371   0.25318077974146663   0.5393377494602607   0.2901912604271057   0.3308554362082618   0.01063526821766662   0.7805303509456989   0.7907756774935695   0.19663847515782248   0.6948919590833847   0.42215247290063596   0.9491896474785065   0.6966937296359754   0.6780052554637713   0.17201305420540866   0.856716158999442   0.8464154257405588   0.4421952614986866   0.7104833320455682   0.09423444156918186   0.062431453488314435   0.11030417972720737   0.7613930513539342   0.4883842440498392   0.37043807986497734   0.8571233999857407   0.22205530189367353   0.19819298362273352   0.03958264365671554   0.8464881317680741   0.44152495094797467   0.40741730612916405   0.8429441684988931   0.15159617268468933   0.019372478047338715
0.4582276586506575   0.14625043886291766   0.473590917220918   0.8473594238419301   0.6015114996512155   0.29983501312235883   0.03139565572223145   0.13687609179636184   0.5072770580820337   0.2374035596340444   0.9210914759950241   0.3754830404424276   0.018892814032194474   0.866965479769067   0.06396807600928336   0.15342773854875405   0.8206998304094609   0.8273828361123515   0.21747994424120928   0.7119027876007794   0.41328252428029694   0.9844386676134584   0.06588377155651995   0.6925303095534407   0.9550548656296394   0.8381882287505408   0.592292854335602   0.8451708857115107   0.3535433659784239   0.538353215628182   0.5608971986133705   0.7082947939151488   0.8462663078963902   0.3009496559941376   0.6398057226183463   0.33281175347272124   0.8273734938641958   0.4339841762250706   0.575837646609063   0.17938401492396716   0.0066736634547348   0.606601340112719   0.35835770236785375   0.46748122732318775   0.5933911391744379   0.6221626724992606   0.29247393081133377   0.774950917769747   0.6383362735447985   0.7839744437487198   0.7001810764757319   0.9297800320582363   0.28479290756637454   0.24562122812053794   0.1392838778623614   0.22148523814308757   0.4385265996699843   0.9446715721264003   0.499478155244015   0.8886734846703663   0.6111531058057885   0.5106873959013298   0.923640508634952   0.7092894697463992
0.6044794423510538   0.9040860557886107   0.5652828062670983   0.24180824242321147   0.011088303176615903   0.28192338328935007   0.27280887545576443   0.4668573246534644   0.37275202963181747   0.4979489395406302   0.5726277989800326   0.5370772925952281   0.08795912206544289   0.25232771142009225   0.43334392111767117   0.31559205445214045   0.6494325223954586   0.3076561392936919   0.9338657658736562   0.4269185697817741   0.03827941658966999   0.7969687433923621   0.010225257238704186   0.717629100035375   0.4337999742386162   0.8928826876037514   0.44494245097160595   0.4758208576121634   0.4227116710620003   0.6109593043144014   0.1721335755158415   0.008963532958699007   0.04995964143018287   0.11301036477377119   0.5995057765358089   0.471886240363471   0.96200051936474   0.860682653353679   0.16616185541813772   0.1562941859113305   0.3125679969692814   0.553026514059987   0.23229608954448153   0.7293756161295564   0.2742885803796114   0.7560577706676249   0.22207083230577734   0.011746516094181526   0.8404886061409952   0.8631750830638736   0.7771283813341714   0.5359256584820181   0.4177769350789949   0.2522157787494722   0.6049948058183299   0.5269621255233191   0.367817293648812   0.139205413975701   0.0054890292825210294   0.05507588515984811   0.40581677428407203   0.2785227606220221   0.8393271738643833   0.8987816992485176
0.09324877731479062   0.725496246562035   0.6070310843199018   0.1694060831189612   0.8189601969351792   0.96943847589441   0.3849602520141244   0.15765956702477965   0.978471590794184   0.10626339283053653   0.607831870679953   0.6217339085427616   0.5606946557151891   0.8540476140810643   0.002837064861623117   0.09477178301944247   0.1928773620663771   0.7148422001053634   0.9973480355791021   0.03969589785959436   0.787060587782305   0.4363194394833413   0.15802086171471877   0.14091419861107676   0.6938118104675145   0.7108231929213062   0.550989777394817   0.9715081154921156   0.8748516135323352   0.7413847170268962   0.16602952538069252   0.8138485484673359   0.8963800227381512   0.6351213241963597   0.5581976547007395   0.1921146399245744   0.33568536702296214   0.7810737101152954   0.5553605898391164   0.0973428569051319   0.14280800495658505   0.066231510009932   0.5580125542600143   0.057646959045537544   0.35574741717428   0.6299120705265907   0.39999169254529554   0.9167327604344607   0.6619356067067655   0.9190888776052845   0.8490019151504785   0.9452246449423451   0.7870839931744302   0.17770416057838823   0.682972389769786   0.13137609647500925   0.890703970436279   0.5425828363820285   0.12477473506904653   0.9392614565504349   0.5550186034133169   0.7615091262667332   0.5694141452299302   0.8419185996453029
0.41221059845673186   0.6952776162568012   0.011401590969915871   0.7842716405997654   0.05646318128245186   0.06536554573021049   0.6114098984246203   0.8675388801653047   0.3945275745756863   0.14627666812492607   0.7624079832741418   0.9223142352229594   0.6074435814012561   0.9685725075465379   0.0794355935043558   0.7909381387479502   0.7167396109649771   0.4259896711645093   0.9546608584353092   0.8516766821975154   0.1617210075516602   0.6644805448977761   0.3852467132053791   0.009758082552212374   0.7495104090949284   0.9692029286409749   0.37384512223546323   0.22548644195244696   0.6930472278124765   0.9038373829107644   0.7624352238108429   0.3579475617871423   0.29851965323679014   0.7575607147858384   0.000027240536701083305   0.43563332656418285   0.6910760718355341   0.7889882072393005   0.9205916470323453   0.6446951878162327   0.974336460870557   0.3629985360747912   0.965930788597036   0.7930185056187173   0.8126154533188968   0.6985179911770151   0.5806840753916569   0.7832604230665049   0.06310504422396848   0.7293150625360402   0.20683895315619363   0.557773981114058   0.370057816411492   0.8254776796252757   0.4444037293453507   0.19982641932691567   0.07153816317470185   0.06791696483943732   0.44437648880864966   0.7641930927627328   0.3804620913391678   0.2789287576001368   0.5237848417763044   0.11949790494650016
0.4061256304686108   0.9159302215253456   0.5578540531792684   0.32647939932778286   0.593510177149714   0.21741223034833052   0.9771699777876115   0.5432189762612779   0.5304051329257454   0.48809716781229034   0.7703310246314179   0.98544499514722   0.16034731651425346   0.6626194881870147   0.3259272952860671   0.7856185758203043   0.0888091533395516   0.5947025233475773   0.8815508064774175   0.02142548305757142   0.7083470620003838   0.31577376574744054   0.35776596470111305   0.9019275781110713   0.30222143153177305   0.39984354422209495   0.7999119115218447   0.5754481787832884   0.7087112543820591   0.18243131387376443   0.8227419337342332   0.03222920252201051   0.17830612145631367   0.694334146061474   0.05241090910281537   0.046784207374790596   0.017958804942060203   0.0317146578744594   0.7264836138167483   0.26116563155448635   0.9291496516025086   0.43701213452688203   0.8449328073393308   0.23974014849691494   0.2208025896021248   0.12123836877944151   0.4871668426382178   0.33781257038584367   0.9185811580703518   0.7213948245573466   0.6872549311163731   0.7623643916025553   0.20986990368829264   0.5389635106835822   0.8645129973821399   0.7301351890805448   0.03156378223197898   0.844629364622108   0.8121020882793245   0.6833509817057541   0.013604977289918779   0.8129147067476487   0.08561847446257623   0.4221853501512678
0.08445532568741017   0.3759025722207666   0.24068566712324538   0.18244520165435288   0.8636527360852854   0.2546642034413251   0.7535188244850276   0.8446326312685092   0.9450715780149337   0.5332693788839785   0.0662638933686545   0.08226823966595394   0.735201674326641   0.9943058682003963   0.20175089598651463   0.35213305058540917   0.703637892094662   0.14967650357828832   0.3896488077071901   0.668782068879655   0.6900329148047433   0.33676179683063967   0.30403033324461387   0.24659671872838718   0.6055775891173331   0.960859224609873   0.06334466612136849   0.0641515170740343   0.7419248530320477   0.7061950211685479   0.30982584163634086   0.21951888580552512   0.796853275017114   0.17292564228456944   0.24356194826768637   0.13725064613957116   0.06165160069047305   0.17861977408417304   0.041811052281171754   0.785117595554162   0.35801370859581105   0.028943270505884695   0.6521622445739816   0.116335526674507   0.6679807937910678   0.6921814736752451   0.34813191132936777   0.8697388079461198   0.06240320467373474   0.731322249065372   0.2847872452079993   0.8055872908720855   0.32047835164168703   0.025127227896824006   0.9749614035716584   0.5860684050665604   0.523625076624573   0.8522015856122546   0.731399455303972   0.4488177589269892   0.4619734759341   0.6735818115280815   0.6895884030228002   0.6637001633728272
0.10395976733828893   0.6446385410221969   0.037426158448818615   0.5473646366983203   0.43597897354722115   0.9524570673469518   0.6892942471194509   0.6776258287522005   0.3735757688734864   0.22113481828157985   0.40450700191145156   0.8720385378801149   0.053097417231799345   0.19600759038475585   0.42954559833979317   0.2859701328135545   0.5294723406072264   0.3438060047725013   0.6981461430358211   0.8371523738865653   0.06749886467312635   0.6702241932444197   0.008557740013020888   0.17345221051373802   0.9635390973348374   0.02558565222222288   0.9711315815642023   0.6260875738154178   0.5275601237876163   0.07312858487527106   0.28183733444475145   0.9484617450632173   0.15398435491412987   0.8519937665936912   0.8773303325332998   0.07642320718310246   0.10088693768233052   0.6559861762089354   0.4477847341935067   0.7904530743695479   0.5714145970751042   0.3121801714364341   0.7496385911576855   0.9533007004829828   0.5039157324019778   0.6419559781920143   0.7410808511446647   0.7798484899692447   0.5403766350671404   0.6163703259697915   0.7699492695804624   0.15376091615382695   0.01281651127952414   0.5432417410945204   0.48811193513571094   0.20529917109060958   0.8588321563653942   0.6912479745008292   0.6107816026024111   0.1288759639075071   0.7579452186830637   0.035261798291893846   0.1629968684089044   0.3384228895379591
0.18653062160795955   0.7230816268554597   0.4133582772512189   0.3851221890549764   0.6826148892059817   0.08112564866344535   0.6722774261065542   0.6052736990857317   0.1422382541388413   0.4647553226936538   0.9023281565260918   0.4515127829319048   0.12942174285931715   0.9215135815991334   0.4142162213903809   0.2462136118412952   0.2705895864939229   0.23026560709830418   0.8034346187879697   0.11733764793378806   0.5126443678108591   0.19500380880641033   0.6404377503790654   0.7789147583958289   0.32611374620289957   0.4719221819509506   0.22707947312784652   0.3937925693408525   0.6434988569969179   0.39079653328750524   0.5548020470212923   0.7885188702551208   0.5012606028580766   0.9260412105938514   0.6524738904952005   0.337006087323216   0.37183885999875943   0.004527628994718013   0.23825766910481963   0.09079247548192083   0.10124927350483653   0.7742620218964138   0.43482305031684987   0.9734548275481327   0.5886049056939774   0.5792582130900035   0.7943852999377845   0.19454006915230385   0.2624911594910778   0.1073360311390529   0.567305826809938   0.8007474998114513   0.6189923024941599   0.7165394978515477   0.012503779788645659   0.012228629556330544   0.11773169963608335   0.7904982872576962   0.36002988929344515   0.6752225422331145   0.7458928396373239   0.7859706582629782   0.12177222018862552   0.5844300667511937
0.6446435661324874   0.011708636366564384   0.6869491698717757   0.610975239203061   0.05603866043850999   0.43245042327656086   0.8925638699339912   0.4164351700507571   0.7935475009474322   0.325114392137508   0.3252580431240532   0.6156876702393057   0.17455519845327228   0.6085748942859603   0.3127542633354075   0.6034590406829752   0.05682349881718892   0.8180766070282641   0.9527243740419624   0.9282364984498607   0.310930659179865   0.03210594876528588   0.8309521538533369   0.343806431698667   0.6662870930473777   0.020397312398721498   0.1440029839815612   0.7328311924956061   0.6102484326088676   0.5879468891221606   0.25143911404757   0.31639602244484905   0.8167009316614354   0.2628324969846526   0.9261810709235169   0.7007083522055433   0.6421457332081631   0.6542576026986923   0.6134268075881093   0.09724931152256812   0.5853222343909743   0.8361809956704281   0.6607024335461469   0.16901281307270746   0.27439157521110924   0.8040750469051423   0.8297502796928101   0.8252063813740405   0.6081044821637316   0.7836777345064209   0.6857472957112489   0.09237518887843438   0.9978560495548641   0.1957308453842602   0.43430818166367885   0.7759791664335853   0.18115511789342859   0.9328983483996076   0.508127110740162   0.07527081422804206   0.5390093846852654   0.2786407457009153   0.8947003031520527   0.9780215027054739
0.9536871502942912   0.4424597500304871   0.2339978696059058   0.8090086896327665   0.679295575083182   0.6383847031253448   0.40424758991309573   0.983802308258726   0.07119109291945028   0.8547069686189239   0.7185002942018468   0.8914271193802916   0.07333504336458625   0.6589761232346637   0.28419211253816795   0.11544795294670629   0.8921799254711577   0.7260777748350562   0.776065001798006   0.04017713871866422   0.3531705407858923   0.4474370291341409   0.8813646986459532   0.062155636013190275   0.3994833904916011   0.004977279103653821   0.6473668290400474   0.2531469463804238   0.7201878154084191   0.366592575978309   0.2431192391269517   0.26934463812169773   0.6489967224889689   0.511885607359385   0.5246189449251049   0.3779175187414061   0.5756616791243827   0.8529094841247213   0.24042683238693688   0.2624695657946998   0.6834817536532249   0.12683170928966517   0.46436183058893094   0.22229242707603558   0.3303112128673327   0.6793946801555243   0.5829971319429778   0.1601367910628453   0.9308278223757316   0.6744174010518704   0.9356303029029304   0.9069898446824215   0.21064000696731244   0.3078248250735614   0.6925110637759787   0.6376452065607238   0.5616432844783436   0.7959392177141763   0.16789211885087382   0.2597276878193177   0.9859816053539608   0.943029733589455   0.927465286463937   0.9972581220246179
0.3024998517007359   0.8161980242997898   0.463103455875006   0.7749656949485824   0.9721886388334032   0.13680334414426554   0.8801063239320283   0.614828903885737   0.04136081645767155   0.4623859430923951   0.9444760210290979   0.7078390592033155   0.8307208094903591   0.15456111801883374   0.2519649572531193   0.0701938526425917   0.26907752501201554   0.35862190030465746   0.08407283840224544   0.810466164823274   0.28309591965805464   0.4155921667152025   0.1566075519383085   0.8132080427986561   0.9805960679573188   0.5993941424154127   0.6935040960633024   0.038242347850073785   0.008407429123915556   0.46259079827114713   0.8133977721312742   0.4234134439643368   0.967046612666244   0.00020485517875203237   0.8689217511021763   0.7155743847610213   0.1363258031758849   0.8456437371599183   0.616956793849057   0.6453805321184296   0.8672482781638694   0.48702183685526085   0.5328839554468116   0.8349143672951556   0.5841523585058147   0.07142967014005837   0.37627640350850305   0.021706324496499448   0.603556290548496   0.4720355277246457   0.6827723074452006   0.9834639766464257   0.5951488614245805   0.009444729453498531   0.8693745353139264   0.5600505326820889   0.6281022487583364   0.009239874274746498   0.0004527842117501477   0.8444761479210676   0.4917764455824515   0.1635961371148282   0.38349599036269316   0.19909561580263807
0.6245281674185821   0.6765743002595673   0.8506120349158816   0.3641812485074825   0.04037580891276741   0.6051446301195089   0.47433563140737856   0.34247492401098306   0.4368195183642714   0.1331091023948633   0.791563323962178   0.3590109473645574   0.841670656939691   0.12366437294136476   0.9221887886482515   0.7989604146824685   0.21356840818135459   0.11442449866661826   0.9217360044365014   0.9544842667614009   0.7217919625989031   0.9508283615517901   0.5382400140738083   0.7553886509587628   0.09726379518032097   0.27425406129222274   0.6876279791579266   0.3912074024512803   0.05688798626755356   0.6691094311727137   0.2132923477505481   0.04873247844029724   0.6200684679032822   0.5360003287778504   0.4217290237883701   0.6897215310757399   0.7783978109635912   0.4123359558364857   0.4995402351401186   0.8907611163932714   0.5648294027822366   0.29791145716986744   0.5778042307036172   0.9362768496318705   0.8430374401833335   0.3470830956180774   0.039564216629808954   0.18088819867310768   0.7457736450030125   0.07282903432585466   0.35193623747188235   0.7896807962218274   0.6888856587354589   0.4037196031531409   0.13864388972133423   0.7409483177815301   0.06881719083217679   0.8677192743752904   0.7169148659329642   0.05122678670579032   0.2904193798685857   0.45538331853880476   0.21737463079284552   0.16046567031251896
0.7255899770863491   0.1574718613689373   0.6395704000892283   0.22418882068064847   0.8825525369030157   0.8103887657508599   0.6000061834594194   0.04330062200754077   0.1367788919000032   0.7375597314250053   0.24806994598753704   0.25361982578571335   0.44789323316454427   0.3338401282718643   0.10942605626620279   0.5126715080041833   0.3790760423323675   0.46612085389657393   0.39251119033323867   0.46144472129839287   0.08865666246378184   0.010737535357769164   0.17513655954039317   0.3009790509858739   0.36306668537743275   0.8532656739888319   0.5355661594511648   0.07679023030522547   0.48051414847441704   0.04287690823797196   0.9355599759917455   0.03348960829768469   0.34373525657441384   0.3053171768129667   0.6874900300042084   0.7798697825119714   0.8958420234098695   0.9714770485411024   0.5780639737380057   0.2671982745077881   0.516765981077502   0.5053561946445284   0.18555278340476694   0.8057535532093952   0.4281093186137202   0.4946186592867593   0.010416223864373783   0.5047745022235213   0.06504263323628748   0.6413529852979274   0.4748500644132089   0.4279842719182958   0.5845284847618705   0.5984760770599554   0.5392900884214634   0.39449466362061114   0.2407932281874566   0.29315890024698876   0.851800058417255   0.6146248811086398   0.34495120477758706   0.32168185170588637   0.27373608467924937   0.3474266066008517
0.828185223700085   0.816325657061358   0.08818330127448243   0.5416730533914564   0.4000759050863648   0.3217069977745986   0.07776707741010866   0.036898551167935195   0.3350332718500773   0.6803540124766712   0.6029170129968997   0.6089142792496394   0.7505047870882069   0.08187793541671573   0.06362692457543626   0.21441961562902825   0.5097115589007503   0.788719035169727   0.21182686615818122   0.5997947345203885   0.16476035412316326   0.4670371834638406   0.9380907814789319   0.2523681279195368   0.33657513042307824   0.6507115264024826   0.8499074802044494   0.7106950745280803   0.9364992253367135   0.32900452862788404   0.7721404027943407   0.6737965233601451   0.6014659534866361   0.6486505161512128   0.16922338979744103   0.06488224411050572   0.8509611663984292   0.5667725807344971   0.10559646522200478   0.8504626284814775   0.34124960749767896   0.7780535455647701   0.8937695990638236   0.250667893961089   0.1764892533745157   0.3110163621009296   0.9556788175848917   0.9982997660415522   0.8399141229514374   0.6603048356984469   0.10577133738044231   0.2876046915134719   0.9034148976147239   0.33130030707056285   0.33363093458610155   0.6138081681533268   0.3019489441280878   0.6826497909193501   0.16440754478866051   0.5489259240428211   0.4509877777296586   0.11587721018485292   0.058811079566655745   0.6984632955613437
0.10973817023197961   0.3378236646200828   0.16504148050283218   0.44779540160025466   0.9332489168574639   0.02680730251915321   0.20936266291794048   0.4494956355587024   0.09333479390602646   0.3665024668207063   0.10359132553749816   0.16189094404523052   0.18991989629130246   0.03520215975014343   0.7699603909513966   0.5480827758919037   0.8879709521632146   0.3525523688307934   0.6055528461627361   0.9991568518490825   0.43698317443355605   0.23667515864594046   0.5467417665960803   0.3006935562877389   0.32724500420157643   0.8988514940258577   0.38170028609324813   0.8528981546874843   0.3939960873441125   0.8720441915067045   0.17233762317530768   0.40340251912878183   0.30066129343808606   0.5055417246859982   0.06874629763780951   0.24151157508355134   0.1107413971467836   0.47033956493585477   0.2987859066864129   0.6934287991916477   0.22277044498356896   0.11778719610506136   0.6932330605236768   0.694271947342565   0.785787270550013   0.8811120374591209   0.14649129392759652   0.3935783910548261   0.4585422663484365   0.9822605434332632   0.7647910078343484   0.5406802363673419   0.06454617900432395   0.1102163519265587   0.5924533846590407   0.13727771723856   0.7638848855662379   0.6046746272405605   0.5237070870212311   0.8957661421550087   0.6531434884194542   0.13433506230470577   0.22492118033481825   0.20233734296336103
0.4303730434358853   0.01654786619964439   0.5316881198111414   0.508065395620796   0.6445857728858724   0.1354358287405235   0.3851968258835449   0.11448700456596983   0.1860435065374359   0.15317528530726032   0.6204058180491966   0.573806768198628   0.12149732753311193   0.04295893338070163   0.027952433390155833   0.43652905096006794   0.3576124419668741   0.43828430614014113   0.5042453463689246   0.5407629088050593   0.7044689535474198   0.30394924383543537   0.27932416603410637   0.33842556584169825   0.2740959101115345   0.287401377635791   0.747636046222965   0.8303601702209022   0.6295101372256622   0.15196554889526748   0.36243922033942005   0.7158731656549325   0.4434666306882262   0.9987902635880072   0.7420334022902235   0.1420663974563045   0.3219693031551143   0.9558313302073055   0.7140809689000677   0.7055373464962366   0.9643568611882403   0.5175470240671644   0.20983562253114305   0.16477443769117725   0.2598879076408204   0.21359778023172904   0.9305114564970367   0.826348871849479   0.9857919975292859   0.926196402595938   0.1828754102740717   0.9959887016285767   0.3562818603036238   0.7742308537006706   0.8204361899346516   0.2801155359736442   0.9128152296153975   0.7754405901126634   0.07840278764442812   0.13804913851733971   0.5908459264602832   0.8196092599053579   0.3643218187443604   0.4325117920211032
0.6264890652720431   0.3020622358381935   0.1544861962132174   0.2677373543299259   0.3666011576312226   0.08846445560646449   0.22397473971618076   0.44138848248044693   0.38080916010193666   0.1622680530105264   0.041099329442109055   0.4453997808518702   0.024527299798312842   0.3880371993098558   0.22066313950745742   0.165284244878226   0.11171207018291528   0.6125966091971924   0.1422603518630293   0.027235106360886288   0.5208661437226321   0.7929873492918345   0.7779385331186688   0.5947233143397831   0.894377078450589   0.49092511345364087   0.6234523369054514   0.3269859600098572   0.5277759208193664   0.4024606578471764   0.3994775971892707   0.8855974775294103   0.14696676071742976   0.24019260483665   0.35837826774716164   0.44019769667754005   0.12243946091911692   0.8521554055267941   0.1377151282397042   0.2749134517993141   0.01072739073620164   0.23955879632960184   0.9954547763766749   0.2476783454384278   0.48986124701356965   0.4465714470377674   0.2175162432580061   0.6529550310986446   0.5954841685629806   0.9556463335841265   0.5940639063525547   0.3259690710887875   0.06770824774361422   0.5531856757369501   0.19458630916328398   0.44037159355937716   0.9207414870261844   0.3129930709003001   0.8362080414161224   0.0001738968818370966   0.7983020261070676   0.46083766537350596   0.6984929131764182   0.7252604450825231
0.7875746353708659   0.2212788690439041   0.7030381367997433   0.47758209964409526   0.29771338835729627   0.7747074220061366   0.4855218935417372   0.8246270685454505   0.7022292197943156   0.8190610884220102   0.8914579871891826   0.4986579974566631   0.6345209720507015   0.26587541268506004   0.6968716780258986   0.05828640389728597   0.7137794850245169   0.95288234178476   0.8606636366097762   0.05811250701544887   0.9154774589174494   0.492044676411254   0.16217072343335798   0.3328520619329258   0.1279028235465835   0.2707658073673499   0.4591325866336147   0.8552699622888306   0.8301894351892872   0.4960583853612132   0.9736106930918775   0.03064289374338   0.12796021539497154   0.6769972969392031   0.08215270590269504   0.5319848962867169   0.49343924334427014   0.41112188425414303   0.3852810278767965   0.4736984923894309   0.7796597583197532   0.45823954246938314   0.5246173912670203   0.415585985373982   0.8641822994023037   0.9661948660581291   0.36244666783366236   0.08273392344105618   0.7362794758557203   0.6954290586907793   0.9033140812000476   0.22746396115222559   0.9060900406664331   0.19937067332956607   0.9297033881081701   0.19682106740884558   0.7781298252714615   0.522373376390363   0.847550682205475   0.6648361711221287   0.2846905819271914   0.11125149213621995   0.46226965432867856   0.19113767873269782
0.5050308236074382   0.6530119496668368   0.9376522630616582   0.7755516933587158   0.6408485242051344   0.6868170836087076   0.5752055952279959   0.6928177699176596   0.9045690483494142   0.9913880249179284   0.6718915140279481   0.46535380876543403   0.9984790076829811   0.7920173515883624   0.742188125919778   0.2685327413565885   0.22034918241151968   0.2696439751979994   0.894637443714303   0.6036965702344598   0.9356586004843284   0.15839248306177942   0.43236778938562437   0.41255889150176195   0.43062777687689013   0.5053805333949426   0.4947155263239662   0.6370071981430462   0.7897792526717557   0.818563449786235   0.9195099310959703   0.9441894282253865   0.8852102043223415   0.8271754248683065   0.24761841706802223   0.47883561945995246   0.8867311966393604   0.0351580732799442   0.5054302911482442   0.21030287810336395   0.6663820142278407   0.7655140980819448   0.6107928474339412   0.6066063078689042   0.7307234137435124   0.6071216150201655   0.17842505804831685   0.19404741636714226   0.3000956368666222   0.10174108162522284   0.6837095317243507   0.5570402182240961   0.5103163841948665   0.2831776318389879   0.7641996006283803   0.6128507899987097   0.625106179872525   0.4560022069706814   0.5165811835603581   0.1340151705387572   0.7383749832331646   0.4208441336907372   0.011150892412113877   0.9237122924353932
0.07199296900532398   0.6553300356087923   0.4003580449781726   0.31710598456648903   0.34126955526181163   0.0482084205886269   0.2219329869298558   0.12305856819934675   0.04117391839518942   0.9464673389634041   0.5382234552055052   0.5660183499752506   0.5308575342003229   0.6632897071244162   0.7740238545771249   0.953167559976541   0.9057513543277979   0.20728750015373476   0.25744267101676677   0.8191523894377838   0.16737637109463324   0.7864433664629976   0.24629177860465293   0.8954400970023906   0.09538340208930926   0.13111333085420526   0.8459337336264803   0.5783341124359016   0.7541138468274976   0.08290491026557835   0.6240007466966244   0.4552755442365548   0.7129399284323082   0.1364375713021743   0.08577729149111933   0.8892571942613042   0.1820823942319853   0.47314786417775817   0.3117534369139945   0.9360896342847632   0.2763310399041874   0.26586036402402335   0.05431076589722768   0.11693724484697939   0.10895466880955415   0.4794169975610258   0.8080189872925747   0.22149714784458882   0.01357126672024489   0.34830366670682056   0.9620852536660944   0.6431630354086872   0.25945741989274723   0.26539875644124217   0.33808450696947   0.18788749117213246   0.546517491460439   0.1289611851390679   0.25230721547835067   0.2986302969108283   0.36443509722845374   0.6558133209613097   0.9405537785643562   0.3625406626260651
0.08810405732426632   0.3899529569372864   0.8862430126671286   0.24560341777908573   0.9791493885147121   0.9105359593762606   0.07822402537455378   0.024106269934496896   0.9655781217944672   0.5622322926694401   0.11613877170845929   0.38094323452580964   0.70612070190172   0.29683353622819786   0.7780542647389893   0.19305574335367715   0.15960321044128098   0.16787235108912998   0.5257470492606386   0.8944254464428488   0.7951681132128272   0.5120590301278202   0.5851932706962824   0.5318847838167837   0.7070640558885609   0.12210607319053383   0.6989502580291539   0.28628136603769805   0.7279146673738488   0.21157011381427324   0.6207262326546   0.2621750961032011   0.7623365455793815   0.6493378211448332   0.5045874609461408   0.8812318615773915   0.05621584367766145   0.3525042849166353   0.7265331962071515   0.6881761182237144   0.8966126332363805   0.18463193382750534   0.2007861469465129   0.7937506717808654   0.10144452002355321   0.6725729036996851   0.6155928762502305   0.2618658879640817   0.3943804641349923   0.5504668305091512   0.9166426182210766   0.9755845219263837   0.6664657967611435   0.33889671669487803   0.2959163855664766   0.7134094258231826   0.904129251181762   0.6895588955500449   0.7913289246203358   0.832177564245791   0.8479134075041006   0.3370546106334095   0.06479572841318433   0.1440014460220767
0.9513007742677201   0.15242267680590418   0.8640095814666714   0.3502507742412112   0.8498562542441669   0.47984977310621907   0.2484167052164409   0.08838488627712948   0.45547579010917466   0.9293829425970678   0.33177408699536426   0.11280036435074578   0.7890099933480311   0.5904862259021898   0.03585770142888763   0.3993909385275632   0.8848807421662691   0.9009273303521449   0.2445287768085518   0.5672133742817721   0.03696733466216846   0.5638727197187353   0.1797330483953675   0.42321192825969545   0.08566656039444832   0.41145004291283116   0.3157234669286961   0.0729611540184842   0.2358103061502814   0.931600269806612   0.06730676171225516   0.9845762677413548   0.7803345160411068   0.002217327209544296   0.7355326747168909   0.871775903390609   0.9913245226930757   0.4117311013073546   0.6996749732880033   0.47238496486304576   0.1064437805268066   0.5108037709552097   0.4551461964794515   0.9051715905812736   0.06947644586463814   0.9469310512364743   0.275413148084084   0.48195966232157816   0.9838098854701898   0.5354810083236432   0.9596896811553879   0.408998508303094   0.7479995793199083   0.6038807385170311   0.8923829194431327   0.4244222405617393   0.9676650632788016   0.6016634113074868   0.15685024472624184   0.5526463371711303   0.976340540585726   0.18993231000013222   0.45717527143823855   0.08026137230808457
0.8698967600589194   0.6791285390449225   0.002029074958787075   0.17508978172681097   0.8004203141942813   0.7321974878084483   0.7266159268747031   0.6931301194052328   0.8166104287240914   0.1967164794848051   0.7669262457193151   0.2841316111021388   0.06861084940418302   0.592835740967774   0.8745433262761824   0.8597093705403995   0.1009457861253814   0.9911723296602872   0.7176930815499405   0.3070630333692692   0.12460524553965542   0.801240019660155   0.26051781011170194   0.22680166106118466   0.25470848548073605   0.12211148061523248   0.2584887351529149   0.05171187933437368   0.4542881712864548   0.38991399280678424   0.5318728082782118   0.3585817599291409   0.6376777425623634   0.19319751332197913   0.7649465625588967   0.07445014882700209   0.5690668931581804   0.6003617723542051   0.8904032362827143   0.21474077828660254   0.46812110703279897   0.6091894426939178   0.1727101547327738   0.9076777449173333   0.34351586149314356   0.8079494230337627   0.9121923446210718   0.6808760838561487   0.0888073760124075   0.6858379424185302   0.653703609468157   0.629164204521775   0.6345192047259527   0.29592394961174606   0.12183080118994515   0.27058244459263414   0.9968414621635893   0.10272643628976692   0.35688423863104846   0.19613229576563204   0.42777456900540894   0.5023646639355618   0.4664810023483342   0.9813915174790295
0.9596534619726099   0.8931752212416441   0.2937708476155604   0.07371377256169616   0.6161376004794664   0.08522579820788126   0.3815785029944886   0.39283768870554747   0.5273302244670589   0.399387855789351   0.7278748935263316   0.7636734841837725   0.8928110197411062   0.10346390617760494   0.6060440923363865   0.49309103959113837   0.895969557577517   0.0007374698878380148   0.249159853705338   0.29695874382550635   0.468194988572108   0.4983728059522762   0.7826788513570038   0.3155672263464768   0.508541526599498   0.6051975847106321   0.48890800374144344   0.24185345378478068   0.8924039261200316   0.5199717865027509   0.10732950074695484   0.8490157650792332   0.36507370165297276   0.12058393071339993   0.3794546072206232   0.08534228089546071   0.4722626819118665   0.017120024535794986   0.7734105148842367   0.5922512413043224   0.5762931243343495   0.016382554647956973   0.5242506611788987   0.29529249747881603   0.10809813576224153   0.5180097486956808   0.7415718098218949   0.9797252711323392   0.5995566091627434   0.9128121639850486   0.25266380608045147   0.7378718173475585   0.7071526830427118   0.3928403774822977   0.14533430533349664   0.8888560522683253   0.3420789813897391   0.2722564467688978   0.7658796981128734   0.8035137713728646   0.8698162994778725   0.25513642223310284   0.9924691832286368   0.21126253006854226
0.29352317514352305   0.23875386758514586   0.46821852204973796   0.9159700325897262   0.18542503938128152   0.7207441188894651   0.726646712227843   0.936244761457387   0.5858684302185381   0.8079319549044164   0.4739829061473916   0.19837294410982853   0.8787157471758262   0.4150915774221187   0.32864860081389496   0.3095168918415032   0.5366367657860871   0.14283513065322087   0.5627689027010215   0.5060031204686386   0.6668204663082146   0.8876987084201181   0.5702997194723849   0.29474059040009637   0.3732972911646915   0.6489448408349722   0.10208119742264686   0.3787705578103701   0.18787225178341   0.9282007219455072   0.37543448519480377   0.4425257963529831   0.602003821564872   0.12026876704109073   0.9014515790474121   0.24415285224315456   0.7232880743890457   0.705177189618972   0.5728029782335172   0.9346359604016513   0.1866513086029586   0.5623420589657512   0.010034075532495655   0.4286328399330127   0.5198308422947441   0.6746433505456331   0.4397343560601108   0.13389224953291634   0.14653355113005254   0.02569850971066088   0.3376531586374639   0.7551216917225462   0.9586612993466426   0.09749778776515372   0.9622186734426602   0.3125958953695631   0.35665747778177054   0.977229020724063   0.06076709439524798   0.06844304312640856   0.6333694033927249   0.27205183110509096   0.4879641161617308   0.13380708272475725
0.4467180947897662   0.7097097721393398   0.4779300406292351   0.7051742427917446   0.9268872524950222   0.03506642159370674   0.03819568456912432   0.5712819932588282   0.7803537013649696   0.00936791188304586   0.7005425259316603   0.816160301536282   0.8216924020183272   0.9118701241178921   0.7383238524890002   0.5035644061667189   0.46503492423655657   0.9346411033938291   0.6775567580937523   0.43512136304031035   0.8316655208438317   0.6625892722887382   0.18959264193202147   0.30131428031555313   0.3849474260540655   0.9528795001493984   0.7116626013027864   0.5961400375238086   0.4580601735590433   0.9178130785556916   0.673466916733662   0.024858044264980367   0.6777064721940737   0.9084451666726457   0.9729243908020017   0.20869774272869834   0.8560140701757465   0.9965750425547536   0.23460053831300143   0.7051333365619794   0.39097914593919   0.061933939160924475   0.5570437802192492   0.27001197352166906   0.5593136250953582   0.39934466687218634   0.36745113828722775   0.968697693206116   0.17436619904129266   0.44646516672278797   0.6557885369844414   0.37255765568230736   0.7163060254822493   0.5286520881670964   0.9823216202507794   0.34769961141732697   0.03859955328817563   0.6202069214944507   0.009397229448777727   0.13900186868862863   0.1825854831124291   0.6236318789396971   0.7747966911357763   0.4338685321266492
0.7916063371732391   0.5616979397787726   0.21775291091652713   0.16385655860498016   0.23229271207788096   0.16235327290658624   0.8503017726292994   0.19515886539886423   0.057926513036588294   0.7158881061837983   0.194513235644858   0.8226012097165569   0.341620487554339   0.1872360180167019   0.21219161539407863   0.4749015982992299   0.30302093426616333   0.5670290965222513   0.20279438594530091   0.33589972961060127   0.12043545115373427   0.9433972175825542   0.4279976948095246   0.902031197483952   0.32882911398049514   0.38169927780378166   0.21024478389299747   0.7381746388789718   0.09653640190261417   0.21934600489719538   0.3599430112636981   0.5430157734801077   0.03860988886602588   0.5034578987133971   0.1654297756188401   0.7204145637635507   0.6969894013116869   0.3162218806966952   0.9532381602247615   0.24551296546432086   0.3939684670455235   0.749192784174444   0.7504437742794605   0.9096132358537196   0.27353301589178924   0.8057955665918898   0.322446079469936   0.007582038369767561   0.9447039019112942   0.4240962887881081   0.11220129557693848   0.2694073994907957   0.8481675000086799   0.2047502838909127   0.7522582843132404   0.7263916260106881   0.8095576111426541   0.7012923851775156   0.5868285086944003   0.005977062247137274   0.11256820983096719   0.38507050448082036   0.6335903484696388   0.7604640967828165
0.7185997427854437   0.6358777203063765   0.8831465741901783   0.8508508609290968   0.4450667268936544   0.8300821537144867   0.5607004947202423   0.8432688225593292   0.5003628249823603   0.40598586492637856   0.44849919914330383   0.5738614230685336   0.6521953249736803   0.20123558103546585   0.6962409148300635   0.8474697970578455   0.8426377138310261   0.4999431958579503   0.10941240613566316   0.8414927348107083   0.730069504000059   0.11487269137712988   0.4758220576660243   0.08102863802789184   0.011469761214615359   0.47899497107075345   0.5926754834758461   0.23017777709879503   0.566403034320961   0.6489128173562668   0.031974988755603784   0.3869089545394658   0.06604020933860072   0.24292695242988824   0.5834757896123   0.8130475314709322   0.41384488436492045   0.0416913713944224   0.8872348747822365   0.9655777344130867   0.5712071705338942   0.5417481755364721   0.7778224686465733   0.12408499960237844   0.8411376665338353   0.4268754841593423   0.30200041098054903   0.04305636157448659   0.8296679053192199   0.9478805130885888   0.7093249275047029   0.8128785844756916   0.2632648709982589   0.29896769573232196   0.6773499387490991   0.4259696299362258   0.19722466165965816   0.056040743302433735   0.0938741491367992   0.6129220984652936   0.7833797772947377   0.01434937190801133   0.2066392743545627   0.6473443640522069
0.21217260676084349   0.4726011963715392   0.42881680570798936   0.5232593644498285   0.3710349402270083   0.04572571221219692   0.12681639472744033   0.48020300287534184   0.5413670349077884   0.09784519912360813   0.4174914672227374   0.6673244183996503   0.2781021639095295   0.7988775033912862   0.7401415284736382   0.2413547884634245   0.08087750224987135   0.7428367600888525   0.6462673793368391   0.628432689998131   0.2974977249551336   0.7284873881808411   0.43962810498227634   0.9810883259459241   0.08532511819429012   0.2558861918093019   0.010811299274287022   0.45782896149609564   0.7142901779672819   0.210160479597105   0.8839949045468467   0.9776259586207537   0.17292314305949344   0.11231528047349684   0.4665034373241093   0.3103015402211035   0.894820979149964   0.3134377770822107   0.7263619088504711   0.06894675175767899   0.8139434769000926   0.5706010169933583   0.08009452951363205   0.44051406175954805   0.5164457519449589   0.8421136288125172   0.6404664245313557   0.45942573581362395   0.43112063375066884   0.5862274370032153   0.6296551252570687   0.0015967743175283413   0.716830455783387   0.3760669574061103   0.745660220710222   0.023970815696774558   0.5439073127238936   0.2637516769326135   0.27915678338611266   0.713669275475671   0.6490863335739296   0.9503138998504028   0.5527948745356416   0.6447225237179921
0.835142856673837   0.3797128828570445   0.4727003450220095   0.20420846195844403   0.31869710472887813   0.5375992540445274   0.8322339204906538   0.74478272614482   0.8875764709782094   0.951371817041312   0.20257879523358516   0.7431859518272917   0.17074601519482233   0.5753048596352017   0.4569185745233632   0.7192151361305171   0.6268387024709288   0.31155318270258825   0.17776179113725055   0.005545860654846092   0.9777523688969991   0.3612392828521855   0.624966916601609   0.36082333693685403   0.1426095122231621   0.981526399995141   0.15226657157959944   0.15661487497841   0.823912407494284   0.44392714595061367   0.32003265108894563   0.41183214883359   0.9363359365160747   0.49255532890930165   0.11745385585536049   0.6686461970062982   0.7655899213212524   0.9172504692740999   0.6605352813319973   0.9494310608757811   0.13875121885032354   0.6056972865715117   0.48277349019474675   0.943885200220935   0.1609988499533244   0.2444580037193262   0.8578065735931378   0.5830618632840809   0.0183893377301623   0.26293160372418517   0.7055400020135384   0.42644698830567096   0.19447693023587834   0.8190044577735714   0.3855073509245927   0.014614839472081023   0.25814099371980365   0.32644912886426986   0.2680534950692322   0.3459686424657828   0.49255107239855134   0.4091986595901699   0.6075182137372349   0.3965375815900017
0.3537998535482278   0.8035013730186582   0.12474472354248817   0.45265238136906666   0.19280100359490338   0.5590433692993321   0.2669381499493504   0.8695905180849857   0.17441166586474108   0.29611176557514685   0.561398147935812   0.4431435297793147   0.9799347356288628   0.47710730780157534   0.17589079701121932   0.4285286903072337   0.7217937419090591   0.15065817893730551   0.9078373019419871   0.08256004784145089   0.22924266951050776   0.7414595193471356   0.30031908820475217   0.6860224662514492   0.87544281596228   0.9379581463284774   0.175574364662264   0.23337008488238256   0.6826418123673766   0.3789147770291454   0.9086362147129137   0.3637795667973969   0.5082301465026355   0.08280301145399856   0.3472380667771016   0.9206360370180822   0.5282954108737727   0.6056957036524232   0.17134726976588227   0.49210734671084855   0.8065016689647136   0.4550375247151177   0.2635099678238952   0.40954729886939767   0.5772589994542059   0.7135780053679821   0.9631908796191431   0.7235248326179484   0.701816183491926   0.7756198590395047   0.787616514956879   0.49015474773556583   0.019174371124549335   0.39670508201035926   0.8789803002439653   0.12637518093816896   0.5109442246219138   0.3139020705563607   0.5317422334668638   0.20573914392008674   0.9826488137481411   0.7082063669039375   0.3603949637009815   0.7136317972092382
0.17614714478342738   0.2531688421888198   0.09688499587708631   0.3040844983398405   0.5988881453292215   0.5395908368208377   0.13369411625794328   0.5805596657218921   0.8970719618372955   0.763970977781333   0.3460776013010643   0.09040491798632624   0.8778975907127462   0.36726589577097385   0.4670973010570989   0.9640297370481573   0.3669533660908324   0.053363825214613116   0.9353550675902351   0.7582905931280706   0.38430455234269134   0.3451574583106756   0.5749601038892537   0.04465879591883238   0.20815740755926393   0.09198861612185581   0.47807510801216735   0.7405742975789918   0.6092692622300424   0.5523977793010181   0.34438099175422404   0.16001463185709974   0.7121973003927469   0.788426801519685   0.9983033904531597   0.0696097138707735   0.8342997096800007   0.4211609057487112   0.5312060893960608   0.1055799768226162   0.46734634358916827   0.36779708053409804   0.5958510218058257   0.34728938369454565   0.08304179124647695   0.02263962222342242   0.0208909179165721   0.3026305877757133   0.874884383687213   0.9306510061015666   0.5428158099044048   0.5620562901967214   0.2656151214571706   0.3782532268005485   0.19843481815018074   0.4020416583396217   0.5534178210644237   0.5898264252808636   0.20013142769702097   0.33243194446884816   0.719118111384423   0.1686655195321524   0.6689253383009601   0.22685196764623197
0.25177176779525473   0.8008684389980544   0.07307431649513438   0.8795625839516863   0.16872997654877778   0.778228816774632   0.05218339857856227   0.5769319961759731   0.29384559286156475   0.8475778106730654   0.5093675886741575   0.014875705979251664   0.028230471404394167   0.4693245838725168   0.3109327705239768   0.61283404763963   0.4748126503399705   0.8794981585916533   0.11080134282695579   0.28040210317078185   0.7556945389555475   0.7108326390595009   0.4418760045259957   0.05355013552454986   0.5039227711602927   0.9099642000614465   0.3688016880308613   0.17398755157286352   0.33519279461151497   0.13173538328681456   0.31661828945229903   0.5970555553968905   0.041347201749950206   0.28415757261374924   0.8072507007781415   0.5821798494176388   0.013116730345556037   0.8148329887412324   0.49631793025416476   0.9693458017780088   0.5383040800055856   0.9353348301495792   0.385516587427209   0.6889436986072269   0.7826095410500381   0.22450219109007838   0.9436405829012133   0.6353935630826771   0.2786867698897454   0.3145379910286319   0.574838894870352   0.4614060115098136   0.9434939752782304   0.18280260774181734   0.258220605418053   0.8643504561129232   0.9021467735282802   0.8986450351280681   0.45096990463991143   0.2821706066952843   0.8890300431827242   0.08381204638683566   0.9546519743857467   0.31282480491727555
0.3507259631771386   0.14847721623725646   0.5691353869585377   0.6238811063100486   0.5681164221271006   0.9239750251471781   0.6254948040573244   0.9884875432273715   0.2894296522373552   0.6094370341185462   0.05065590918697237   0.5270815317175579   0.34593567695912475   0.4266344263767289   0.7924353037689194   0.6627310756046348   0.4437889034308445   0.5279893912486607   0.341465399129008   0.38056046890935047   0.5547588602481204   0.4441773448618251   0.3868134247432613   0.06773566399207491   0.2040328970709817   0.2957001286245686   0.8176780377847236   0.4438545576820263   0.6359164749438811   0.3717251034773906   0.1921832337273992   0.45536701445465483   0.34648682270652603   0.7622880693588443   0.14152732454042685   0.9282854827370969   0.0005511457474013225   0.3356536429821155   0.34909202077150747   0.2655544071324621   0.5567622423165568   0.8076642517334547   0.007626621642499515   0.8849939382231117   0.0020033820684364836   0.36348690687162966   0.6208131968992382   0.8172582742310367   0.7979704849974548   0.06778677824706102   0.8031351591145146   0.3734037165490104   0.1620540100535736   0.6960616747696705   0.6109519253871154   0.9180367020943556   0.8155671873470476   0.9337736054108261   0.4694246008466886   0.9897512193572587   0.8150160415996462   0.5981199624287107   0.1203325800751811   0.7241968122247966
0.2582537992830894   0.7904557106952559   0.1127059584326816   0.839202874001685   0.2562504172146529   0.4269688038236263   0.49189276153344336   0.021944599770648297   0.45827993221719815   0.35918202557656526   0.6887576024189287   0.6485408832216378   0.29622592216362453   0.6631203508068948   0.07780567703181329   0.7305041811272823   0.480658734816577   0.7293467453960687   0.6083810761851247   0.7407529617700236   0.6656426932169308   0.13122678296735804   0.4880484961099436   0.016556149545226904   0.4073888939338414   0.3407710722721021   0.375342537677262   0.17735327554354188   0.1511384767191885   0.9138022684484759   0.8834497761438187   0.15540867577289358   0.6928585445019904   0.5546202428719106   0.19469217372488995   0.5068677925512557   0.3966326223383658   0.8914998920650158   0.11688649669307664   0.7763636114239735   0.9159738875217888   0.16215314666894717   0.5085054205079519   0.035610649653949895   0.25033119430485795   0.030926363701589125   0.02045692439800833   0.019054500108722987   0.8429423003710166   0.690155291429487   0.6451143867207463   0.8417012245651811   0.691803823651828   0.7763530229810112   0.7616646105769277   0.6862925487922875   0.9989452791498377   0.2217327801091005   0.5669724368520377   0.1794247562410318   0.6023126568114718   0.3302328880440847   0.4500859401589611   0.40306114481705835
0.6863387692896831   0.1680797413751375   0.9415805196510092   0.36745049516310846   0.43600757498482506   0.13715337767354838   0.9211235952530008   0.34839599505438545   0.5930652746138085   0.4469980862440614   0.2760092085322545   0.5066947704892044   0.9012614509619805   0.6706450632630503   0.5143445979553268   0.8204022216969169   0.9023161718121429   0.44891228315394976   0.9473721611032891   0.6409774654558851   0.300003515000671   0.1186793951098651   0.497286220944328   0.2379163206388267   0.6136647457109881   0.9505996537347275   0.5557057012933189   0.8704658254757183   0.17765717072616297   0.8134462760611793   0.6345821060403181   0.5220698304213328   0.5845918961123544   0.3664481898171178   0.35857289750806354   0.015375059932128394   0.683330445150374   0.6958031265540675   0.8442282995527367   0.19497283823521153   0.7810142733382311   0.24689084340011777   0.8968561384494476   0.5539953727793264   0.4810107583375601   0.12821144829025266   0.3995699175051196   0.31607905214049975   0.8673460126265721   0.17761179455552506   0.8438642162118007   0.4456132266647815   0.6896888419004091   0.36416551849434586   0.20928211017148265   0.9235433962434487   0.10509694578805465   0.9977173286772281   0.8507092126634191   0.9081683363113203   0.4217665006376807   0.3019142021231605   0.006480913110682403   0.7131954980761088
0.6407522272994496   0.05502335872304273   0.1096247746612348   0.15920012529678235   0.15974146896188948   0.9268119104327901   0.7100548571561152   0.8431210731562826   0.29239545633531744   0.749200115877265   0.8661906409443145   0.3975078464915011   0.6027066144349084   0.3850345973829191   0.6569085307728318   0.4739644502480524   0.4976096686468537   0.3873172687056911   0.8061993181094127   0.565796113936732   0.07584316800917298   0.08540306658253058   0.7997184049987303   0.8526006158606233   0.43509094070972343   0.030379707859487844   0.6900936303374955   0.6934004905638409   0.2753494717478339   0.10356779742669778   0.9800387731813803   0.8502794174075583   0.9829540154125165   0.35436768154943277   0.11384813223706582   0.4527715709160572   0.3802474009776082   0.9693330841665136   0.456939601464234   0.9788071206680048   0.8826377323307545   0.5820158154608226   0.6507402833548213   0.4130110067312727   0.8067945643215815   0.496612748878292   0.851021878356091   0.5604103908706495   0.3717036236118581   0.46623304101880414   0.16092824801859545   0.8670099003068086   0.0963541518640242   0.3626652435921064   0.18088947483721515   0.016730482899250235   0.11340013645150772   0.008297562042673592   0.06704134260014934   0.563958911983193   0.7331527354738996   0.038964477876159934   0.6101017411359153   0.5851517913151882
0.8505150031431451   0.4569486624153374   0.959361457781094   0.17214078458391555   0.043720438821563526   0.9603359135370454   0.10833957942500311   0.6117303937132661   0.6720168152097055   0.4941028725182412   0.9474113314064077   0.7447204934064575   0.5756626633456812   0.13143762892613484   0.7665218565691925   0.7279900105072074   0.4622625268941735   0.12314006688346124   0.6994805139690432   0.1640310985240143   0.729109791420274   0.08417558900730131   0.08937877283312783   0.578879307208826   0.8785947882771289   0.627226926591964   0.13001731505203376   0.40673852262491045   0.8348743494555654   0.6668910130549186   0.02167773562703066   0.7950081289116444   0.16285753424585997   0.17278814053667738   0.07426640422062301   0.05028763550518679   0.5871948709001787   0.041350511610542526   0.3077445476514305   0.3222976249979795   0.12493234400600524   0.9182104447270812   0.6082640336823874   0.15826652647396516   0.3958225525857313   0.83403485571978   0.5188852608492595   0.5793872192651391   0.5172277643086024   0.20680792912781604   0.3888679457972257   0.1726486966402287   0.682353414853037   0.5399169160728975   0.3671902101701951   0.37764056772858434   0.5194958806071771   0.3671287755362201   0.29292380594957207   0.32735293222339756   0.9323010097069984   0.32577826392567755   0.9851792582981416   0.005055307225418086
0.8073686657009931   0.4075678191985963   0.3769152246157542   0.8467887807514529   0.4115461131152618   0.5735329634788163   0.8580299637664948   0.2674015614863138   0.8943183488066594   0.3667250343510003   0.469162017969269   0.09475286484608507   0.21196493395362237   0.8268081182781029   0.1019718077990739   0.7171122971175007   0.6924690533464453   0.4596793427418827   0.8090480018495019   0.3897593648941032   0.760168043639447   0.13390107881620517   0.8238687435513603   0.3847040576686851   0.9527993779384539   0.7263332596176089   0.44695351893560603   0.5379152769172322   0.5412532648231921   0.1528002961387926   0.5889235551691113   0.27051371543091846   0.6469349160165327   0.7860752617877923   0.1197615371998423   0.17576085058483337   0.4349699820629104   0.9592671435096894   0.0177897294007684   0.45864855346733263   0.7425009287164651   0.49958780076780673   0.20874172755126658   0.06888918857322944   0.9823328850770181   0.36568672195160157   0.3848729839999063   0.6841851309045444   0.029533507138564164   0.6393534623339927   0.9379194650643002   0.14626985398731215   0.48828024231537204   0.48655316619520006   0.34899590989518897   0.8757561385563937   0.8413453262988393   0.7004779044074078   0.2292343726953467   0.6999952879715604   0.4063753442359289   0.7412107608977183   0.2114446432945783   0.24134673450422772
0.6638744155194639   0.24162296012991158   0.002702915743311724   0.1724575459309983   0.6815415304424458   0.87593623817831   0.6178299317434054   0.48827241502645397   0.6520080233038816   0.23658277584431736   0.6799104666791052   0.3420025610391418   0.1637277809885096   0.7500296096491172   0.3309145567839161   0.46624642248274806   0.3223824546896703   0.04955170524170947   0.10168018408856945   0.7662511345111878   0.9160071104537414   0.3083409443439912   0.8902355407939911   0.52490440000696   0.2521326949342775   0.06671798421407958   0.8875326250506794   0.3524468540759617   0.5705911644918317   0.19078174603576956   0.26970269330727403   0.8641744390495077   0.91858314118795   0.9541989701914522   0.5897922266281689   0.522171878010366   0.7548553601994404   0.20416936054233495   0.25887766984425276   0.0559254555276179   0.43247290550977013   0.1546176553006255   0.1571974857556833   0.2896743210164302   0.5164657950560287   0.8462767109566344   0.2669619449616922   0.7647699210094702   0.2643331001217513   0.7795587267425548   0.37942931991101275   0.4123230669335085   0.6937419356299196   0.5887769807067852   0.10972662660373872   0.5481486278840008   0.7751587944419696   0.6345780105153329   0.5199343999755698   0.025976749873634745   0.020303434242529107   0.430408649972998   0.2610567301313171   0.9700512943460169
0.587830528732759   0.2757909946723725   0.10385924437563378   0.6803769733295867   0.07136473367673017   0.4295142837157382   0.8368972994139416   0.9156070523201165   0.8070316335549789   0.6499555569731834   0.4574679795029289   0.503283985386608   0.11328969792505927   0.061178576266398305   0.34774135289919017   0.9551353575026073   0.3381309034830897   0.42660056575106536   0.8278069529236204   0.9291586076289725   0.3178274692405606   0.9961919157780673   0.5667502227923032   0.9591073132829557   0.7299969405078016   0.7204009211056949   0.4628909784166695   0.27873033995336904   0.6586322068310715   0.2908866373899567   0.6259936790027278   0.3631232876332525   0.8516005732760926   0.6409310804167732   0.16852569949979895   0.8598393022466445   0.7383108753510333   0.5797525041503749   0.8207843466006087   0.9047039447440373   0.4001799718679436   0.15315193839930955   0.9929773936769885   0.9755453371150647   0.08235250262738299   0.15696002262124217   0.42622717088468515   0.01643802383210904   0.3523555621195813   0.43655910151554733   0.9633361924680156   0.73770768387874   0.6937233552885098   0.14567246412559065   0.33734251346528776   0.3745843962454875   0.8421227820124172   0.5047413837088174   0.1688168139654888   0.5147450939988429   0.10381190666138393   0.9249888795584426   0.34803246736488   0.6100411492548057
0.7036319347934403   0.7718369411591329   0.35505507368789163   0.6344958121397409   0.6212794321660573   0.6148769185378908   0.9288279028032065   0.6180577883076319   0.268923870046476   0.17831781702234348   0.9654917103351909   0.8803501044288919   0.5752005147579662   0.03264535289675285   0.6281491968699031   0.5057657081834044   0.7330777327455489   0.5279039691879354   0.45933238290441425   0.9910206141845614   0.629265826084165   0.6029150896294929   0.1112999155395342   0.3809794649297558   0.9256338912907247   0.8310781484703599   0.7562448418516425   0.7464836527900148   0.30435445912466735   0.2162012299324691   0.827416939048436   0.1284258644823829   0.03543058907819133   0.0378834129101256   0.8619252287132452   0.24807576005349102   0.46023007432022517   0.005238060013372756   0.23377603184334214   0.7423100518700866   0.7271523415746762   0.4773340908254374   0.7744436489389279   0.7512894376855251   0.09788651549051124   0.8744190011959445   0.6631437333993937   0.3703099727557694   0.17225262419978657   0.04334085272558458   0.9068988915477512   0.6238263199657545   0.8678981650751192   0.8271396227931155   0.0794819524993151   0.4954004554833716   0.8324675759969279   0.7892562098829898   0.21755672378606988   0.24732469542988056   0.3722375016767027   0.7840181498696172   0.9837806919427278   0.505014643559794
0.6450851601020265   0.3066840590441798   0.20933704300379982   0.7537252058742688   0.5471986446115152   0.4322650578482353   0.5461933096044062   0.38341523311849945   0.3749460204117287   0.38892420512265075   0.639294418056655   0.7595889131527449   0.5070478553366095   0.5617845823295352   0.5598124655573399   0.2641884576693733   0.6745802793396816   0.7725283724465454   0.34225574177127   0.016863762239492767   0.30234277766297885   0.9885102225769282   0.3584750498285422   0.5118491186796988   0.6572576175609524   0.6818261635327485   0.14913800682474243   0.75812391280543   0.11005897294943709   0.24956110568451315   0.6029446972203363   0.37470867968693056   0.7351129525377084   0.8606369005618624   0.9636502791636814   0.6151197665341857   0.22806509720109888   0.29885231823232716   0.4038378136063415   0.3509313088648123   0.5534848178614173   0.5263239457857818   0.061582071835071556   0.3340675466253195   0.25114204019843844   0.5378137232088536   0.7031070220065293   0.8222184279456207   0.5938844226374861   0.8559875596761051   0.5539690151817869   0.0640945151401907   0.48382544968804897   0.606426453991592   0.9510243179614506   0.6893858354532602   0.7487124971503406   0.7457895534297295   0.9873740387977692   0.0742660689190745   0.5206473999492417   0.4469372351974024   0.5835362251914277   0.7233347600542622
0.9671625820878245   0.9206132894116206   0.5219541533563561   0.38926721342894266   0.716020541889386   0.382799566202767   0.8188471313498268   0.5670487854833219   0.12213611925189989   0.5268120065266619   0.2648781161680399   0.5029542703431312   0.6383106695638509   0.9203855525350699   0.3138537982065894   0.8135684348898711   0.8895981724135102   0.1745959991053404   0.3264797594088202   0.7393023659707966   0.3689507724642686   0.727658763907938   0.7429435342173926   0.01596760591653441   0.4017881903764442   0.8070454744963174   0.22098938086103645   0.6267003924875917   0.6857676484870582   0.4242459082935504   0.4021422495112097   0.05965160700426977   0.5636315292351584   0.8974339017668884   0.13726413334316978   0.5566973366611385   0.9253208596713074   0.9770483492318185   0.8234103351365805   0.7431289017712673   0.035722687257797134   0.8024523501264781   0.4969305757277602   0.0038265358004707663   0.6667719147935286   0.07479358621854013   0.7539870415103677   0.9878589298839363   0.2649837244170844   0.26774811172222274   0.5329976606493312   0.3611585373963446   0.5792160759300262   0.8435022034286723   0.13085541113812155   0.3015069303920749   0.015584546694867845   0.9460683016617839   0.9935912777949518   0.7448095937309364   0.09026368702356043   0.9690199524299653   0.17018094265837133   0.0016806919596689624
0.05454099976576329   0.1665676023034872   0.6732503669306111   0.9978541561591981   0.3877690849722347   0.09177401608494706   0.9192633254202434   0.009995226275261839   0.12278536055515037   0.8240259043627244   0.3862656647709122   0.6488366888789172   0.5435692846251242   0.9805237009340521   0.25541025363279063   0.3473297584868424   0.5279847379302564   0.03445539927226817   0.2618189758378388   0.602520164755906   0.43772105090669594   0.06543544684230285   0.09163803317946749   0.6008394727962371   0.3831800511409327   0.8988678445388156   0.4183876662488564   0.6029853166370388   0.995410966168698   0.8070938284538686   0.499124340828613   0.592990090361777   0.8726256056135475   0.9830679240911442   0.11285867605770085   0.9441534014828598   0.3290563209884233   0.002544223157092209   0.8574484224249103   0.5968236429960174   0.801071583058167   0.9680888238848241   0.5956294465870714   0.9943034782401114   0.363350532151471   0.9026533770425212   0.5039914134076039   0.3934640054438744   0.9801704810105384   0.003785532503705549   0.08560374715874752   0.7904786888068355   0.9847595148418404   0.19669170404983696   0.5864794063301345   0.1974885984450585   0.11213390922829293   0.21362377995869272   0.4736207302724337   0.2533351969621987   0.7830775882398696   0.21107955680160054   0.6161723078475234   0.6565115539661812
0.9820060051817027   0.24299073291677648   0.020542861260452   0.6622080757260699   0.6186554730302316   0.3403373558742553   0.5165514478528481   0.26874407028219544   0.6384849920196932   0.33655182337054973   0.43094770069410054   0.47826538147535996   0.6537254771778528   0.13986011932071277   0.8444682943639661   0.28077678303030146   0.5415915679495599   0.92623633936202   0.37084756409153236   0.027441586068102743   0.7585139797096903   0.7151567825604195   0.754675256244009   0.3709300321019215   0.7765079745279876   0.472166049643643   0.734132394983557   0.7087219563758517   0.157852501497756   0.13182869376938774   0.21758094713070888   0.4399778860936562   0.5193675094780628   0.795276870398838   0.7866332464366084   0.9617125046182963   0.86564203230021   0.6554167510781252   0.9421649520726423   0.6809357215879948   0.32405046435065016   0.7291804117161051   0.5713173879811099   0.6534941355198921   0.56553648464096   0.01402362915568567   0.816642131737101   0.28256410341797056   0.7890285101129723   0.5418575795120426   0.08250973675354398   0.5738421470421189   0.6311760086152163   0.4100288857426549   0.864928789622835   0.13386426094846274   0.11180849913715353   0.614752015343817   0.07829554318622675   0.1721517563301665   0.24616646683694354   0.9593352642656917   0.13613059111358447   0.4912160347421717
0.9221160024862934   0.2301548525495865   0.5648132031324745   0.8377218992222796   0.3565795178453335   0.21613122339390084   0.7481710713953736   0.555157795804309   0.5675510077323612   0.6742736438818582   0.6656613346418296   0.9813156487621901   0.936374999117145   0.2642447581392033   0.8007325450189946   0.8474513878137274   0.8245664999799914   0.6494927427953864   0.7224370018327678   0.6752996314835609   0.5784000331430479   0.6901574785296947   0.5863064107191833   0.18408359674138922   0.6562840306567544   0.46000262598010816   0.0214932075867088   0.34636169751910956   0.29970451281142096   0.24387140258620732   0.27332213619133516   0.7912039017148005   0.7321535050790597   0.5695977587043491   0.6076608015495055   0.8098882529526104   0.7957785059619149   0.30535300056514586   0.8069282565305109   0.962436865138883   0.9712120059819235   0.6558602577697594   0.08449125469774316   0.2871372336553221   0.39281197283887564   0.9657027792400648   0.49818484397855983   0.10305363691393293   0.7365279421821211   0.5057001532599567   0.476691636391851   0.7566919393948234   0.43682342937070023   0.26182875067374933   0.20336950020051583   0.9654880376800228   0.7046699242916404   0.6922309919694002   0.5957086986510103   0.15559978472741243   0.9088914183297256   0.3868779914042544   0.7887804421204994   0.19316291958852938
0.937679412347802   0.7310177336344948   0.7042891874227561   0.9060256859332073   0.5448674395089265   0.7653149543944301   0.20610434344419634   0.8029720490192743   0.8083394973268052   0.25961480113447344   0.7294127070523453   0.04628010962445098   0.37151606795610503   0.9977860504607241   0.5260432068518295   0.08079207194442815   0.6668461436644646   0.30555505849132397   0.9303345082008192   0.9251922872170157   0.757954725334739   0.9186770670870695   0.14155406608031992   0.7320293676284864   0.8202753129869369   0.18765933345257468   0.43726487865756375   0.826003681695279   0.2754078734780104   0.4223443790581446   0.2311605352133674   0.02303163267600475   0.4670683761512051   0.16272957792367113   0.501747828161022   0.9767515230515538   0.0955523081951001   0.16494352746294696   0.9757046213091926   0.8959594511071256   0.42870616453063554   0.859388468971623   0.04537011310837332   0.9707671638901099   0.6707514391958965   0.9407114018845535   0.9038160470280534   0.23873779626162356   0.8504761262089597   0.7530520684319788   0.46655116837048966   0.41273411456634446   0.5750682527309493   0.33070768937383416   0.23539063315712222   0.38970248189033974   0.10799987657974419   0.16797811145016303   0.7336428049961001   0.41295095883878596   0.012447568384644083   0.003034583987216064   0.7579381836869076   0.5169915077316604
0.5837414038540085   0.14364611501559305   0.7125680705785343   0.5462243438415505   0.912989964658112   0.20293471313103958   0.8087520235504809   0.3074865475799269   0.06251383844915225   0.4498826446990608   0.34220085517999127   0.8947524330135824   0.4874455857182029   0.11917495532522666   0.10681022202286902   0.5050499511232427   0.3794457091384587   0.9511968438750636   0.37316741702676887   0.09209899228445671   0.36699814075381465   0.9481622598878475   0.6152292333398612   0.5751074845527964   0.7832567368998061   0.8045161448722545   0.9026611627613269   0.028883140711245932   0.8702667722416941   0.6015814317412149   0.09390913921084604   0.7213965931313191   0.8077529337925419   0.15169878704215412   0.7517082840308548   0.8266441601177367   0.32030734807433897   0.03252383171692744   0.6448980620079857   0.321594208994494   0.9408616389358803   0.08132698784186382   0.2717306449812169   0.22949521671003725   0.5738634981820656   0.13316472795401624   0.6565014116413557   0.6543877321572409   0.7906067612822595   0.3286485830817617   0.7538402488800288   0.6255045914459949   0.9203399890405654   0.7270671513405468   0.6599311096691827   0.9041079983146759   0.11258705524802345   0.5753683642983927   0.9082228256383279   0.07746383819693925   0.7922797071736845   0.5428445325814653   0.2633247636303422   0.7558696292024453
0.8514180682378042   0.46151754473960144   0.9915941186491253   0.526374412492408   0.27755457005573864   0.3283528167855852   0.3350927070077696   0.8719866803351671   0.48694780877347915   0.9997042337038234   0.5812524581277408   0.24648208888917225   0.5666078197329137   0.27263708236327666   0.9213213484585582   0.34237409057449636   0.4540207644848903   0.697268718064884   0.013098522820230262   0.2649102523775571   0.6617410573112059   0.15442418548341874   0.7497737591898881   0.5090406231751118   0.8103229890734016   0.6929066407438174   0.7581796405407628   0.9826662106827038   0.532768419017663   0.36455382395823216   0.42308693353299326   0.11067953034753658   0.0458206102441839   0.36484959025440866   0.8418344754052524   0.8641974414583643   0.47921279051127014   0.09221250789113201   0.9205131269466942   0.521823350883868   0.02519202602637979   0.394943789826248   0.9074146041264639   0.2569130985063109   0.3634509687151739   0.24051960434282926   0.15764084493657585   0.747872475331199   0.5531279796417723   0.5476129635990119   0.399461204395813   0.7652062646484953   0.020359560624109256   0.1830591396407798   0.9763742708628197   0.6545267343009588   0.9745389503799253   0.8182095493863711   0.13453979545756736   0.7903292928425943   0.49532615986865525   0.7259970414952391   0.21402666851087315   0.2685059419587264
0.4701341338422754   0.33105325166899113   0.30661206438440924   0.011592843452415513   0.10668316512710152   0.09053364732616184   0.1489712194478334   0.26372036812121646   0.5535551854853292   0.5429206837271499   0.7495100150520204   0.4985141034727211   0.53319562486122   0.35986154408637006   0.7731357441892006   0.8439873691717624   0.5586566744812946   0.5416519946999989   0.6385959487316333   0.05365807632916806   0.06333051461263939   0.8156549532047598   0.4245692802207601   0.7851521343704416   0.593196380770364   0.4846017015357687   0.1179572158363509   0.7735592909180261   0.48651321564326244   0.3940680542096069   0.9689859963885175   0.5098389227968098   0.9329580301579332   0.851147370482457   0.21947598133649712   0.011324819324088556   0.3997624052967132   0.4912858263960869   0.4463402371472965   0.16733745015232612   0.8411057308154186   0.949633831696088   0.8077442884156631   0.11367937382315807   0.7777752162027792   0.1339788784913281   0.3831750081949031   0.3285272394527164   0.18457883543241524   0.6493771769555594   0.2652177923585522   0.5549679485346902   0.6980656197891528   0.2553091227459525   0.2962317959700347   0.045129025737880545   0.7651075896312196   0.40416175226349554   0.07675581463353758   0.03380420641379199   0.3653451843345064   0.9128759258674086   0.6304155774862411   0.8664667562614659
0.5242394535190879   0.9632420941713207   0.822671289070578   0.7527873824383078   0.7464642373163086   0.8292632156799925   0.4394962808756748   0.4242601429855914   0.5618854018838935   0.17988603872443312   0.17427848851712266   0.8692921944509011   0.8638197820947406   0.9245769159784806   0.878046692547088   0.8241631687130206   0.09871219246352099   0.5204151637149851   0.8012908779135504   0.7903589622992286   0.7333670081290146   0.6075392378475765   0.1708753004273093   0.9238922060377628   0.2091275546099267   0.6442971436762558   0.3482040113567314   0.17110482359945495   0.4626633172936181   0.8150339279962633   0.9087077304810566   0.7468446806138636   0.9007779154097246   0.6351478892718302   0.7344292419639339   0.8775524861629624   0.03695813331498404   0.7105709732933495   0.8563825494168459   0.05338931744994179   0.9382459408514631   0.19015580957836448   0.05509167150329551   0.26303035515071316   0.2048789327224485   0.582616571730788   0.8842163710759862   0.3391381491129504   0.9957513781125218   0.9383194280545322   0.5360123597192549   0.16803332551349545   0.5330880608189037   0.12328550005826887   0.6273046292381983   0.4211886448996319   0.6323101454091791   0.4881376107864387   0.8928753872742644   0.5436361587366695   0.595352012094195   0.7775666374930892   0.03649283785741849   0.49024684128672774
0.6571060712427319   0.5874108279147247   0.981401166354123   0.22721648613601456   0.45222713852028346   0.004794256183936702   0.09718479527813677   0.8880783370230642   0.45647576040776167   0.06647482812940454   0.561172435558882   0.7200450115095687   0.923387699588858   0.9431893280711356   0.9338678063206837   0.29885636660993675   0.2910775541796789   0.45505171728469695   0.04099241904641923   0.7552202078732673   0.6957255420854839   0.6774850797916078   0.004499581189000741   0.2649733665865395   0.038619470842751975   0.09007425187688312   0.023098414834877765   0.03775688045052497   0.5863923323224686   0.0852799956929464   0.925913619556741   0.14967854342746084   0.12991657191470685   0.018805167563541874   0.3647411839978591   0.42963353191789216   0.20652887232584888   0.07561583949240622   0.43087337767717543   0.1307771653079554   0.91545131814617   0.6205641222077093   0.3898809586307562   0.37555695743468814   0.21972577606068602   0.9430790424161014   0.3853813774417555   0.11058359084814863   0.18110630521793405   0.8530047905392183   0.3622829626068777   0.07282671039762366   0.5947139728954656   0.7677247948462719   0.4363693430501367   0.9231481669701628   0.46479740098075867   0.7489196272827301   0.07162815905227762   0.49351463505227067   0.2582685286549098   0.6733037877903238   0.6407547813751022   0.36273746974431526
0.34281721050873987   0.05273966558261458   0.250873822744346   0.9871805123096271   0.1230914344480538   0.10966062316651314   0.8654924453025905   0.8765969214614785   0.9419851292301198   0.2566558326272948   0.5032094826957129   0.8037702110638548   0.3472711563346542   0.48893103778102287   0.06684013964557611   0.8806220440936919   0.8824737553538955   0.7400114104982929   0.9952119805932985   0.3871074090414213   0.6242052266989857   0.066707622707969   0.3544571992181963   0.024369939297106052   0.2813880161902459   0.013967957125354417   0.10358337647385032   0.03718942698747896   0.15829658174219208   0.9043073339588413   0.23809093117125982   0.1605925055260005   0.21631145251207234   0.6476515013315465   0.734881448475547   0.3568222944621457   0.8690402961774181   0.1587204635505236   0.6680413088299709   0.4762002503684537   0.9865665408235226   0.4187090530522308   0.6728293282366724   0.08909284132703241   0.36236131412453687   0.3520014303442618   0.3183721290184761   0.06472290202992635   0.08097329793429096   0.33803347321890737   0.21478875254462576   0.027533475042447405   0.9226767161920989   0.4337261392600661   0.9766978213733659   0.866940969516447   0.7063652636800265   0.7860746379285196   0.24181637289781896   0.5101186750543012   0.8373249675026084   0.627354174377996   0.5737750640678481   0.0339184246858475
0.8507584266790859   0.2086451213257652   0.9009457358311757   0.9448255833588151   0.488397112554549   0.8566436909815034   0.5825736068126995   0.8801026813288887   0.407423814620258   0.5186102177625961   0.36778485426807384   0.8525692062864413   0.48474709842815916   0.08488407850253002   0.39108703289470786   0.9856282367699944   0.7783818347481326   0.29880944057401043   0.14927065999688893   0.4755095617156932   0.9410568672455242   0.6714552661960145   0.5754955959290409   0.4415911370298457   0.09029844056643832   0.46281014487024924   0.6745498600978652   0.4967655536710306   0.6019013280118893   0.6061664538887458   0.09197625328516557   0.6166628723421419   0.1944775133916313   0.08755623612614971   0.7241913990170917   0.7640936660557005   0.7097304149634722   0.0026721576236196963   0.33310436612238387   0.7784654292857062   0.9313485802153396   0.7038627170496092   0.18383370612549493   0.3029558675700129   0.9902917129698154   0.03240745085359481   0.6083381101964541   0.8613647305401673   0.8999932724033771   0.5695973059833456   0.9337882500985889   0.3645991768691366   0.2980919443914878   0.9634308520945998   0.8418119968134233   0.7479363045269948   0.10361443099985647   0.8758746159684501   0.11762059779633162   0.9838426384712943   0.3938840160363843   0.8732024583448303   0.7845162316739478   0.2053772091855881
0.46253543582104467   0.16933974129522109   0.6006825255484528   0.9024213416155752   0.4722437228512293   0.13693229044162628   0.9923444153519987   0.04105661107540795   0.5722504504478522   0.5673349844582807   0.058556165253409787   0.6764574342062714   0.2741585060563644   0.6039041323636809   0.21674416843998642   0.9285211296792766   0.1705440750565079   0.728029516395231   0.0991235706436548   0.9446784912079823   0.7766600590201236   0.8548270580504005   0.31460733896970705   0.7393012820223942   0.3141246231990789   0.6854873167551795   0.7139248134212542   0.836879940406819   0.8418809003478497   0.5485550263135531   0.7215803980692556   0.7958233293314111   0.2696304498999975   0.9812200418552725   0.6630242328158458   0.11936589512513979   0.9954719438436331   0.3773159094915915   0.4462800643758593   0.1908447654458632   0.8249278687871252   0.6492863930963606   0.3471564937322045   0.24616627423788087   0.04826780976700161   0.7944593350459601   0.03254915476249743   0.5068649922154866   0.7341431865679227   0.10897201829078063   0.3186243413412432   0.6699850518086675   0.892262286220073   0.5604169919772275   0.5970439432719877   0.8741617224772564   0.6226318363200755   0.579196950121955   0.934019710456142   0.7547958273521167   0.6271598924764423   0.2018810406303635   0.48773964608028264   0.5639510619062534
0.8022320236893171   0.5525946475340029   0.14058315234807817   0.3177847876683726   0.7539642139223155   0.7581353124880428   0.10803399758558073   0.810919795452886   0.01982102735439284   0.6491632941972622   0.7894096562443376   0.1409347436442184   0.1275587411343198   0.08874630222003473   0.19236571297234986   0.266773021166962   0.5049269048142443   0.5095493520980797   0.25834600251620793   0.5119771938148453   0.877767012337802   0.3076683114677162   0.7706063564359252   0.9480261319085919   0.0755349886484848   0.7550736639337133   0.6300232040878471   0.6302413442402193   0.3215707747261693   0.9969383514456706   0.5219892065022663   0.8193215487873333   0.30174974737177646   0.3477750572484083   0.7325795502579289   0.6783868051431149   0.17419100623745662   0.2590287550283736   0.5402138372855789   0.41161378397615295   0.6692641014232124   0.7494794029302939   0.28186783476937105   0.8996365901613076   0.7914970890854104   0.44181109146257763   0.5112614783334458   0.9516104582527157   0.7159621004369255   0.6867374275288644   0.8812382742455988   0.3213691140124964   0.3943913257107563   0.6897990760831938   0.3592490677433324   0.502047565225163   0.09264157833897985   0.3420240188347855   0.6266695174854036   0.8236607600820481   0.9184505721015233   0.08299526380641192   0.08645568019982458   0.4120469761058952
0.24918647067831093   0.33351586087611806   0.8045878454304536   0.5124103859445875   0.45768938159290057   0.8917047694135404   0.29332636709700777   0.5607999276918718   0.741727281155975   0.2049673418846761   0.41208809285140907   0.23943081367937535   0.3473359554452187   0.5151682658014822   0.0528390251080767   0.7373832484542123   0.2546943771062389   0.17314424696669678   0.42616950762267314   0.9137224883721642   0.3362438050047156   0.09014898316028484   0.33971382742284856   0.5016755122662689   0.08705733432640471   0.7566331222841668   0.535125981992395   0.9892651263216815   0.6293679527335041   0.8649283528706264   0.2417996148953873   0.4284651986298097   0.8876406715775291   0.6599610109859503   0.8297115220439782   0.18903438495043434   0.5403047161323105   0.144792745184468   0.7768724969359015   0.45165113649622207   0.2856103390260716   0.9716484982177712   0.3507029893132284   0.5379286481240579   0.949366534021356   0.8814995150574864   0.0109891618903798   0.03625313585778893   0.8623091996949512   0.1248663927733196   0.47586317989798477   0.046988009536107475   0.2329412469614471   0.2599380399026932   0.23406356500259745   0.6185228109062978   0.34530057538391795   0.599977028916743   0.4043520429586192   0.42948842595586345   0.8049958592516075   0.455184283732275   0.6274795460227176   0.9778372894596414
0.519385520225536   0.4835357855145037   0.27677655670948925   0.4399086413355835   0.57001898620418   0.6020362704570174   0.26578739481910946   0.40365550547779455   0.7077097865092287   0.4771698776836978   0.7899242149211247   0.3566674959416871   0.47476853954778164   0.21723183778100455   0.5558606499185272   0.7381446850353893   0.12946796416386366   0.6172548088642615   0.15150860695990806   0.3086562590795258   0.3244721049122562   0.16207052513198664   0.5240290609371904   0.33081896961988444   0.8050865846867202   0.6785347396174829   0.24725250422770115   0.890910328284301   0.2350675984825403   0.07649846916046553   0.9814651094085917   0.48725482280650634   0.5273578119733116   0.5993285914767678   0.19154089448746697   0.13058732686481925   0.05258927242552997   0.38209675369576324   0.6356802445689397   0.39244264182942995   0.9231213082616663   0.7648419448315016   0.48417163760903165   0.0837863827499041   0.5986492033494101   0.602771419699515   0.9601425766718412   0.7529674131300197   0.7935626186626898   0.9242366800820321   0.71289007244414   0.8620570848457187   0.5584950201801495   0.8477382109215665   0.7314249630355484   0.3748022620392124   0.03113720820683797   0.2484096194447988   0.5398840685480815   0.24421493517439313   0.9785479357813079   0.8663128657490357   0.9042038239791418   0.8517722933449632
0.0554266275196417   0.10147092091753399   0.4200321863701101   0.767985910595059   0.4567774241702316   0.498699501218019   0.45988960969826886   0.015018497465039395   0.6632148055075417   0.5744628211359869   0.7469995372541287   0.15296141261932064   0.10471978532739215   0.7267246102144204   0.015574574218580335   0.7781591505801083   0.07358257712055419   0.47831499076962153   0.47569050567049886   0.5339442154057151   0.09503464133924619   0.6120021250205859   0.5714866816913572   0.682171922060752   0.03960801381960449   0.5105312041030519   0.15145449532124705   0.9141860114656929   0.582830589649373   0.011831702885032911   0.6915648856229782   0.8991675140006535   0.9196157841418312   0.43736888174904603   0.9445653483688494   0.7462061013813328   0.8148959988144391   0.7106442715346257   0.9289907741502691   0.9680469508012246   0.7413134216938848   0.23232928076500417   0.45330026847977023   0.4341027353955094   0.6462787803546387   0.6203271557444183   0.881813586788413   0.7519308133347575   0.6066707665350342   0.10979595164136637   0.730359091467166   0.8377448018690646   0.023840176885661254   0.09796424875633346   0.03879420584418782   0.9385772878684111   0.10422439274383004   0.6605953670072875   0.09422885747533837   0.1923711864870783   0.28932839392939097   0.9499510954726618   0.16523808332506926   0.22432423568585372
0.5480149722355061   0.7176218147076576   0.711937814845299   0.7902215002903443   0.9017361918808674   0.0972946589632393   0.8301242280568859   0.03829068695558678   0.2950654253458333   0.987498707321873   0.09976513658971989   0.20054588508652219   0.27122524846017204   0.8895344585655395   0.060970930745532066   0.26196859721811105   0.167000855716342   0.22893909155825204   0.9667420732701937   0.06959741073103276   0.877672461786951   0.2789879960855903   0.8015039899451245   0.8452731750451791   0.32965748955144486   0.5613661813779327   0.08956617509982544   0.05505167475483477   0.4279212976705774   0.4640715224146934   0.25944194704293955   0.01676098779924799   0.13285587232474413   0.47657281509282046   0.15967681045321963   0.8162151027127258   0.8616306238645721   0.587038356527281   0.09870587970768757   0.5542465054946147   0.6946297681482302   0.35809926496902894   0.13196380643749386   0.484649094763582   0.8169573063612792   0.0791112688834387   0.33045981649236944   0.6393759197184029   0.4872998168098343   0.517745087505506   0.240893641392544   0.5843242449635682   0.05937851913925688   0.05367356509081261   0.9814516943496044   0.5675632571643202   0.9265226468145128   0.5771007499979921   0.8217748838963849   0.7513481544515944   0.06489202294994063   0.9900623934707111   0.7230690041886972   0.1971016489569796
0.3702622548017105   0.6319631285016822   0.5911051977512034   0.7124525541933976   0.5533049484404313   0.5528518596182435   0.26064538125883396   0.07307663447499466   0.06600513163059707   0.03510677211273749   0.01975173986629   0.48875238951142647   0.006626612491340191   0.9814332070219248   0.03830004551668554   0.9211891323471063   0.08010396567682744   0.4043324570239327   0.21652516162030072   0.16984097789551192   0.015211942726886809   0.4142700635532216   0.4934561574316034   0.9727393289385323   0.6449496879251763   0.7823069350515394   0.9023509596804   0.2602867747451347   0.09164473948474494   0.2294550754332959   0.6417055784215661   0.18721014027014005   0.02563960785414788   0.19434830332055844   0.6219538385552761   0.6984577507587135   0.019012995362807688   0.21291509629863356   0.5836537930385906   0.7772686184116073   0.9389090296859802   0.8085826392747009   0.36712863141828983   0.6074276405160953   0.9236970869590935   0.3943125757214792   0.8736724739866863   0.6346883115775631   0.27874739903391715   0.6120056406699398   0.9713215143062863   0.3744015368324284   0.18710265954917218   0.3825505652366439   0.3296159358847202   0.18719139656228834   0.1614630516950243   0.18820226191608547   0.7076620973294442   0.48873364580357476   0.1424500563322166   0.9752871656174519   0.1240083042908536   0.7114650273919675
0.20354102664623638   0.1667045263427511   0.7568796728725637   0.10403738687587212   0.27984393968714294   0.7723919506212719   0.8832071988858774   0.46934907529830905   0.0010965406532258094   0.16038630995133205   0.9118856845795911   0.09494753846588067   0.8139938811040536   0.7778357447146882   0.5822697486948708   0.9077561419035923   0.6525308294090293   0.5896334827986027   0.8746076513654267   0.4190224961000175   0.5100807730768127   0.6143463171811507   0.7505993470745731   0.70755746870805   0.30653974643057635   0.44764179083839967   0.9937196742020094   0.6035200818321779   0.026695806743433394   0.6752498402171279   0.11051247531613194   0.13417100653386885   0.025599266090207583   0.5148635302657958   0.19862679073654088   0.03922346806798819   0.21160538498615394   0.7370277855511076   0.6163570420416701   0.13146732616439588   0.5590745555771246   0.1473943027525049   0.7417493906762433   0.7124448300643783   0.04899378250031192   0.5330479855713541   0.9911500436016702   0.004887361356328314   0.7424540360697356   0.08540619473295442   0.997430369399661   0.4013672795241504   0.7157582293263022   0.4101563545158266   0.8869178940835291   0.26719627299028154   0.6901589632360946   0.8952928242500309   0.6882911033469882   0.22797280492229335   0.47855357824994066   0.15826503869892328   0.07193406130531811   0.09650547875789749
0.919479022672816   0.010870735946418396   0.33018467062907475   0.38406064869351914   0.8704852401725041   0.4778227503750643   0.33903462702740444   0.3791732873371908   0.1280312041027685   0.39241655564210987   0.3416042576277435   0.9778060078130404   0.4122729747764663   0.9822602011262832   0.4546863635442145   0.7106097348227589   0.7221140115403717   0.08696737687625238   0.7663952601972264   0.48263692990046553   0.24356043329043103   0.9287023381773291   0.6944611988919082   0.386131451142568   0.324081410617615   0.9178316022309106   0.36427652826283347   0.0020708024490488737   0.4535961704451109   0.4400088518558464   0.02524190123542901   0.6228975151118581   0.3255649663423424   0.047592296213736535   0.6836376436076855   0.6450915072988176   0.913291991565876   0.0653320950874533   0.22895128006347104   0.9344817724760588   0.19117798002550437   0.978364718211201   0.4625560198662447   0.45184484257559326   0.9476175467350734   0.04966238003387184   0.7680948209743365   0.06571339143302524   0.6235361361174584   0.13183077780296115   0.40381829271150305   0.06364258898397637   0.16993996567234745   0.6918219259471148   0.378576391476074   0.4407450738721183   0.844374999330005   0.6442296297333782   0.6949387478683885   0.7956535665733007   0.931083007764129   0.578897534645925   0.46598746780491745   0.861171794097242
0.7399050277386247   0.600532816434724   0.0034314479386727535   0.40932695152164866   0.7922874810035513   0.5508704364008522   0.23533662696433624   0.3436135600886234   0.16875134488609292   0.419039658597891   0.8315183342528332   0.2799709711046471   0.9988113792137455   0.7272177326507763   0.4529419427767592   0.8392258972325287   0.15443637988374037   0.08298810291739804   0.7580031949083706   0.04357233065922805   0.22335337211961137   0.5040905682714731   0.2920157271034532   0.1824005365619861   0.4834483443809867   0.9035577518367491   0.2885842791647804   0.7730735850403374   0.6911608633774354   0.352687315435897   0.05324765220044418   0.429460024951714   0.5224095184913425   0.933647656838006   0.22172931794761097   0.14948905384706693   0.523598139277597   0.20642992418722972   0.7687873751708518   0.3102631566145382   0.3691617593938567   0.12344182126983168   0.010784180262481154   0.26669082595531013   0.1458083872742453   0.6193512529983586   0.7187684531590279   0.08429028939332403   0.6623600428932586   0.7157935011616094   0.4301841739942476   0.3112167043529866   0.9711991795158231   0.36310618572571246   0.3769365217938034   0.8817566794012726   0.4487896610244806   0.42945852888770647   0.15520720384619238   0.7322676255542057   0.9251915217468835   0.22302860470047678   0.3864198286753406   0.4220044689396675
0.5560297623530268   0.0995867834306451   0.37563564841285946   0.15531364298435735   0.4102213750787815   0.48023553043228656   0.6568671952538314   0.0710233535910333   0.747861332185523   0.7644420292706771   0.2266830212595839   0.7598066492380467   0.7766621526696998   0.40133584354496465   0.8497464994657805   0.8780499698367741   0.32787249164521926   0.9718773146572581   0.6945392956195882   0.14578234428256845   0.40268096989833574   0.7488487099567814   0.3081194669442475   0.723777875342901   0.846651207545309   0.6492619265261362   0.9324838185313881   0.5684642323585436   0.43642983246652745   0.16902639609384976   0.27561662327755665   0.49744087876751036   0.6885685002810045   0.40458436682317267   0.048933602017972755   0.7376342295294637   0.9119063476113047   0.003248523278207999   0.1991871025521922   0.8595842596926895   0.5840338559660855   0.031371208620949845   0.5046478069326041   0.7138019154101211   0.18135288606774969   0.28252249866416845   0.19652833998835653   0.9900240400672201   0.33470167852244076   0.6332605721380322   0.26404452145696844   0.42155980770867646   0.8982718460559133   0.46423417604418243   0.9884278981794118   0.9241189289411661   0.2097033457749088   0.059649809221009785   0.939494296161439   0.18648469941170248   0.2977969981636041   0.056401285942801783   0.7403071936092468   0.32690043971901295
0.7137631421975187   0.02503007732185194   0.2356593866766427   0.6130985243088919   0.532410256129769   0.7425075786576835   0.03913104668828616   0.6230744842416718   0.19770857760732827   0.1092470065196513   0.7750865252313177   0.20151467653299537   0.299436731551415   0.6450128304754689   0.7866586270519059   0.2773957475918293   0.08973338577650619   0.585363021254459   0.8471643308904669   0.09091104818012682   0.7919363876129021   0.5289617353116574   0.10685713728122015   0.7640106084611139   0.07817324541538341   0.5039316579898053   0.8711977506045775   0.15091208415222196   0.5457629892856144   0.7614240793321219   0.8320667039162913   0.5278375999105501   0.34805441167828616   0.6521770728124706   0.056980178684973556   0.32632292337755475   0.04861768012687118   0.00716424233700172   0.2703215516330676   0.04892717578572547   0.958884294350365   0.42180122108254264   0.42315722074260065   0.9580161276055986   0.1669479067374629   0.8928394857708853   0.3163000834613805   0.1940055191444848   0.08877466132207948   0.38890782778107996   0.44510233285680306   0.04309343499226283   0.543011672036465   0.627483748448958   0.6130356289405118   0.5152558350817127   0.19495726035817892   0.9753066756364874   0.5560554502555382   0.18893291170415794   0.14633958023130775   0.9681424332994858   0.2857338986224706   0.14000573591843246
0.18745528588094276   0.5463412122169431   0.8625766778798699   0.1819896083128338   0.020507379143479856   0.6535017264460578   0.5462765944184894   0.987984089168349   0.9317327178214003   0.26459389866497784   0.10117426156168641   0.9448906541760862   0.3887210457849353   0.6371101502160198   0.48813863262117463   0.4296348190943735   0.1937637854267564   0.6618034745795324   0.9320831823656365   0.24070190739021557   0.04742420519544866   0.6936610412800466   0.6463492837431658   0.10069617147178313   0.8599689193145059   0.14731982906310345   0.7837726058632959   0.9187065631589493   0.839461540171026   0.4938181026170457   0.23749601144480642   0.9307224739906003   0.9077288223496257   0.2292242039520678   0.13632174988312   0.9858318198145141   0.5190077765646903   0.5921140537360481   0.6481831172619453   0.5561970007201406   0.32524399113793395   0.9303105791565157   0.716099934896309   0.315495093329925   0.2778197859424853   0.23664953787646914   0.0697506511531431   0.21479892185814187   0.4178508666279794   0.08932970881336569   0.2859780452898472   0.29609235869919254   0.5783893264569534   0.59551160619632   0.048482033845040795   0.3653698847085923   0.6706605041073277   0.3662874022442522   0.9121602839619207   0.37953806489407815   0.1516527275426373   0.7741733485082042   0.2639771666999754   0.8233410641739376
0.8264087364047034   0.8438627693516885   0.5478772318036664   0.5078459708440126   0.548588950462218   0.6072132314752193   0.4781265806505233   0.2930470489858707   0.13073808383423863   0.5178835226618537   0.19214853536067614   0.9969546902866782   0.5523487573772853   0.9223719164655336   0.14366650151563534   0.6315848055780859   0.8816882532699576   0.5560845142212814   0.23150621755371456   0.25204674068400773   0.7300355257273203   0.7819111657130772   0.9675290508537392   0.4287056765100702   0.903626789322617   0.9380483963613887   0.4196518190500727   0.9208597056660576   0.3550378388603989   0.3308351648861694   0.9415252383995494   0.6278126566801869   0.22429975502616026   0.8129516422243157   0.7493767030388733   0.6308579663935088   0.671950997648875   0.8905797257587821   0.605710201523238   0.9992731608154228   0.7902627443789174   0.3344952115375007   0.37420398396952337   0.7472264201314152   0.060227218651597074   0.5525840458244236   0.4066749331157842   0.31852074362134497   0.15660042932898013   0.6145356494630348   0.9870231140657114   0.39766103795528734   0.8015625904685812   0.2837004845768654   0.045497875666162084   0.7698483812751005   0.577262835442421   0.4707488423525497   0.2961211726272888   0.13899041488159172   0.905311837793546   0.5801691165937676   0.6904109711040509   0.13971725406616886
0.11504909341462864   0.24567390505626682   0.31620698713452755   0.39249083393475376   0.05482187476303157   0.6930898592318433   0.9095320540187434   0.0739700903134088   0.8982214454340515   0.07855420976880846   0.922508939953032   0.6763090523581214   0.0966588549654702   0.794853725191943   0.8770110642868698   0.906460671083021   0.5193960195230493   0.3241048828393933   0.580889891659581   0.7674702562014293   0.6140841817295032   0.7439357662456257   0.8904789205555301   0.6277530021352604   0.4990350883148746   0.4982618611893589   0.5742719334210025   0.23526216820050663   0.444213213551843   0.8051720019575156   0.6647398794022591   0.16129207788709785   0.5459917681177916   0.7266177921887071   0.7422309394492271   0.4849830255289764   0.4493329131523214   0.9317640669967642   0.8652198751623573   0.5785223544459555   0.9299368936292721   0.6076591841573709   0.28432998350277633   0.8110520982445262   0.31585271189976893   0.863723417911745   0.39385106294724626   0.18329909610926573   0.8168176235848944   0.36546155672238617   0.8195791295262438   0.948036927908759   0.37260441003305134   0.5602895547648705   0.1548392501239846   0.7867448500216613   0.8266126419152597   0.8336717625761634   0.41260831067475745   0.30176182449268485   0.3772797287629384   0.9019076955793993   0.5473884355124001   0.7232394700467295
0.44734283513366624   0.29424851142202846   0.26305845200962374   0.9121873718022033   0.1314901232338973   0.4305250935102834   0.8692073890623775   0.7288882756929376   0.31467249964900296   0.06506353678789725   0.049628259536133756   0.7808513477841785   0.9420680896159516   0.5047739820230267   0.8947890094121491   0.9941064977625172   0.11545544770069184   0.6711022194468633   0.4821806987373917   0.6923446732698324   0.7381757189377535   0.769194523867464   0.9347922632249916   0.9691052032231029   0.2908328838040872   0.4749460124454356   0.6717338112153678   0.05691783142089961   0.1593427605701899   0.0444209189351522   0.8025264221529903   0.32802955572796205   0.8446702609211869   0.979357382147255   0.7528981626168566   0.5471782079437836   0.9026021713052353   0.4745834001242282   0.8581091532047075   0.5530717101812663   0.7871467236045435   0.803481180677365   0.37592845446731576   0.8607270369114339   0.048971004666790025   0.03428665680990085   0.44113619124232417   0.891621833688331   0.7581381208627028   0.5593406443644653   0.7694023800269563   0.8347040022674314   0.5987953602925129   0.5149197254293131   0.966875957873966   0.5066744465394694   0.754125099371326   0.5355623432820581   0.21397779525710936   0.9594962385956858   0.8515229280660906   0.060978943157829854   0.35586864205240193   0.4064245284144195
0.06437620446154718   0.25749776248046496   0.9799401875850862   0.5456974915029855   0.015405199794757154   0.2232111056705641   0.538803996342762   0.6540756578146545   0.25726707893205436   0.6638704613060988   0.7694016163158057   0.8193716555472231   0.6584717186395415   0.14895073587678578   0.8025256584418398   0.3126972090077538   0.9043466192682155   0.6133883925947277   0.5885478631847303   0.35320097041206794   0.05282369120212476   0.5524094494368978   0.23267922113232842   0.9467764419976484   0.9884474867405776   0.2949116869564329   0.2527390335472423   0.4010789504946629   0.9730422869458204   0.0717005812858688   0.7139350372044803   0.7470032926800083   0.715775208013766   0.40783011997977   0.9445334208886746   0.9276316371327852   0.05730348937422468   0.25887938410298417   0.1420077624468349   0.6149344281250314   0.15295687010600925   0.6454909915082565   0.5534598992621046   0.26173345771296347   0.1001331789038845   0.09308154207135862   0.3207806781297761   0.31495701571531504   0.11168569216330691   0.7981698551149258   0.06804164458253385   0.9138780652206522   0.1386434052174865   0.7264692738290569   0.35410660737805355   0.16687477254064376   0.42286819720372043   0.318639153849287   0.40957318648937896   0.23924313540785855   0.36556470782949574   0.059759769746302795   0.267565424042544   0.6243087072828271
0.21260783772348646   0.4142687782380463   0.7141055247804394   0.3625752495698636   0.11247465881960197   0.3211872361666877   0.3933248466506633   0.047618233854548574   0.0007889666562950566   0.523017381051762   0.3252832020681295   0.13374016863389646   0.8621455614388086   0.7965481072227051   0.9711765946900759   0.9668653960932527   0.4392773642350882   0.4779089533734181   0.561603408200697   0.7276222606853942   0.07371265640559244   0.41814918362711534   0.29403798415815297   0.10331355340256704   0.861104818682106   0.003880405389068981   0.5799324593777135   0.7407383038327034   0.748630159862504   0.6826931692223813   0.18660761272705018   0.6931200699781549   0.7478411932062089   0.15967578817061928   0.8613244106589207   0.5593799013442584   0.8856956317674004   0.3631276809479142   0.8901478159688447   0.5925145052510057   0.44641826753231223   0.8852187275744962   0.32854440776814775   0.8648922445656116   0.3727056111267198   0.4670695439473808   0.03450642360999481   0.7615786911630446   0.5116007924446139   0.46318913855831184   0.4545739642322813   0.020840387330341135   0.7629706325821098   0.7804959693359306   0.2679663515052311   0.32772031735218626   0.015129439375900902   0.6208201811653112   0.40664194084631045   0.7683404160079279   0.12943380760850054   0.25769250021739704   0.5164941248774657   0.17582591075692214
0.6830155400761884   0.37247377264290094   0.18794971710931793   0.3109336661913105   0.3103099289494685   0.9054042286955202   0.15344329349932312   0.549354975028266   0.7987091365048548   0.44221509013720833   0.6988693292670418   0.5285145876979248   0.03573850392274489   0.6617191208012778   0.43090297776181063   0.20079427034573857   0.020609064546843987   0.04089893963596651   0.0242610369155002   0.4324538543378107   0.8911752569383434   0.7832064394185695   0.5077669120380345   0.2566279435808886   0.20815971686215512   0.41073266677566855   0.3198171949287166   0.945694277389578   0.8978497879126865   0.5053284380801484   0.16637390142939346   0.39633930236131204   0.09914065140783186   0.06311334794294009   0.46750457216235164   0.8678247146633872   0.06340214748508698   0.4013942271416623   0.036601594400541   0.6670304443176486   0.042793082938242986   0.3604952875056958   0.012340557485040798   0.2345765899798379   0.15161782599989954   0.5772888480871263   0.5045736454470063   0.9779486463989494   0.9434581091377444   0.16655618131145777   0.1847564505182897   0.03225436900937134   0.04560832122505782   0.6612277432313094   0.018382549088896256   0.6359150666480593   0.946467669817226   0.5981143952883693   0.5508779769265446   0.7680903519846721   0.883065522332139   0.196720168146707   0.5142763825260036   0.10105990766702352
0.840272439393896   0.8362248806410112   0.5019358250409628   0.8664833176871856   0.6886546133939965   0.25893603255388487   0.9973621795939565   0.8885346712882363   0.7451965042562521   0.09237985124242709   0.8126057290756667   0.8562803022788649   0.6995881830311943   0.4311521080111177   0.7942231799867705   0.2203652356308056   0.7531205132139683   0.8330377127227484   0.24334520306022595   0.45227488364613344   0.8700549908818292   0.6363175445760414   0.7290688205342223   0.35121497597910994   0.0297825514879333   0.8000926639350302   0.22713299549325952   0.4847316582919243   0.3411279380939368   0.5411566313811453   0.22977081589930304   0.5961969870036881   0.5959314338376848   0.44877678013871825   0.41716508682363623   0.7399166847248232   0.8963432508064905   0.017624672127600518   0.6229419068368657   0.5195514490940176   0.14322273759252221   0.18458695940485212   0.3795967037766398   0.06727656544788416   0.27316774671069294   0.5482694148288108   0.6505278832424174   0.7160615894687742   0.24338519522275961   0.7481767508937806   0.4233948877491579   0.23132993117684988   0.9022572571288228   0.2070201195126352   0.19362407184985486   0.6351329441731618   0.30632582329113806   0.758243339373917   0.7764589850262187   0.8952162594483386   0.40998257248464753   0.7406186672463164   0.15351707818935292   0.375664810354321
0.2667598348921253   0.5560317078414643   0.7739203744127131   0.30838824490643685   0.9935920881814324   0.007762293012653621   0.12339249117029573   0.5923266554376626   0.7502068929586727   0.25958554211887314   0.6999976034211378   0.36099672426081275   0.84794963582985   0.052565422606237935   0.506373531571283   0.725863780087651   0.541623812538712   0.29432208323232095   0.7299145465450643   0.8306475206393124   0.13164124005406438   0.5537034159860046   0.5763974683557114   0.4549827102849914   0.8648814051619391   0.9976717081445402   0.8024770939429983   0.14659446537855453   0.8712893169805067   0.9899094151318866   0.6790846027727024   0.5542678099408919   0.121082424021834   0.7303238730130135   0.9790869993515646   0.19327108568007914   0.27313278819198406   0.6777584504067755   0.4727134677802817   0.4674073055924282   0.7315089756532721   0.38343636717445456   0.7427989212352174   0.6367597849531158   0.5998677355992078   0.82973295118845   0.16640145287950606   0.18177707466812446   0.7349863304372687   0.8320612430439098   0.3639243589365078   0.035182609289569934   0.863697013456762   0.8421518279120233   0.6848397561638053   0.48091479934867803   0.742614589434928   0.11182795489900973   0.7057527568122407   0.28764371366859887   0.46948180124294386   0.4340695044922342   0.23303928903195895   0.8202364080761707
0.7379728255896717   0.05063313731777964   0.4902403677967415   0.18347662312305488   0.13810508999046398   0.22090018612932963   0.3238389149172355   0.0016995484549304134   0.4031187595531953   0.38883894308541983   0.9599145559807276   0.9665169391653605   0.5394217460964333   0.5466871151733966   0.2750747998169223   0.48560213981668243   0.7968071566615055   0.43485916027438687   0.5693220430046817   0.19795842614808357   0.32732535541856156   0.0007896557821526545   0.3362827539727227   0.37772201807191286   0.5893525298288899   0.950156518464373   0.8460423861759812   0.19424539494885798   0.45124743983842586   0.7292563323350434   0.5222034712587457   0.19254584649392756   0.048128680285230534   0.34041738924962356   0.562288915278018   0.2260289073285671   0.5087069341887972   0.793730274076227   0.28721411546109576   0.7404267675118846   0.7118997775272917   0.3588711138018401   0.7178920724564142   0.5424683413638011   0.38457442210873016   0.3580814580196875   0.3816093184836914   0.16474632329188824   0.7952218922798404   0.40792493955531445   0.5355669323077102   0.9705009283430303   0.34397445244141456   0.6786686072202711   0.013363461048964506   0.7779550818491027   0.295845772156184   0.3382512179706475   0.4510745457709464   0.5519261745205356   0.7871388379673868   0.5445209438944205   0.16386043030985067   0.811499407008651
0.07523906044009511   0.18564983009258038   0.4459683578534365   0.26903106564484985   0.6906646383313649   0.8275683720728929   0.06435903936974513   0.10428474235296162   0.8954427460515245   0.41964343251757846   0.5287921070620349   0.13378381400993136   0.55146829361011   0.7409748252973074   0.5154286460130704   0.35582873216082866   0.255622521453926   0.4027236073266599   0.06435410024212397   0.8039025576402931   0.4684836834865391   0.8582026634322394   0.9004936699322733   0.9924031506316422   0.39324462304644403   0.672552833339659   0.45452531207883673   0.7233720849867923   0.7025799847150791   0.8449844612667661   0.39016627270909165   0.6190873426338307   0.8071372386635546   0.42534102874918767   0.8613741656470567   0.48530352862389936   0.25566894505344456   0.6843662034518803   0.34594551963398634   0.12947479646307064   0.00004642359951857744   0.2816425961252204   0.2815914193918624   0.3255722388227775   0.5315627401129794   0.423439932692981   0.3810977494595891   0.3331690881911354   0.1383181170665354   0.750887099353322   0.9265724373807523   0.609797003204343   0.4357381323514563   0.9059026380865559   0.5364061646716607   0.9907096605705124   0.6286008936879017   0.48056160933736825   0.675031999024604   0.505406131946613   0.37293194863445717   0.7961954058854879   0.32908647939061764   0.37593133548354235
0.3728855250349386   0.5145528097602675   0.04749505999875526   0.0503590966607648   0.8413227849219591   0.0911128770672865   0.6663973105391662   0.7171900084696294   0.7030046678554237   0.3402257777139645   0.7398248731584138   0.10739300526528639   0.26726653550396745   0.4343231396274086   0.2034187084867532   0.11668334469477405   0.6386656418160658   0.9537615302900404   0.5283867094621493   0.611277212748161   0.26573369318160855   0.15756612440455248   0.19930023007153164   0.2353458772646187   0.89284816814667   0.6430133146442849   0.15180517007277639   0.1849867806038539   0.051525383224710834   0.5519004375769985   0.4854078595336102   0.4677967721342245   0.3485207153692871   0.21167465986303394   0.7455829863751963   0.3604037668689381   0.08125417986531965   0.7773515202356254   0.5421642778884431   0.24372042217416404   0.4425885380492539   0.823589989945585   0.013777568426293837   0.632443209426003   0.17685484486764536   0.6660238655410324   0.8144773383547622   0.39709733216138426   0.28400667672097535   0.023010550896747507   0.6626721682819858   0.2121105515575304   0.23248129349626453   0.47111011331974906   0.17726430874837562   0.7443137794233059   0.8839605781269775   0.2594354534567151   0.43168132237317935   0.38391001255436785   0.8027063982616578   0.4820839332210898   0.8895170444847362   0.1401895903802038
0.3601178602124039   0.6584939432755048   0.8757394760584424   0.5077463809542008   0.18326301534475853   0.9924700777344724   0.0612621377036802   0.11064904879281653   0.8992563386237832   0.9694595268377248   0.3985899694216944   0.8985384972352861   0.6667750451275186   0.4983494135179758   0.22132566067331874   0.15422471781198024   0.7828144670005412   0.2389139600612607   0.7896443383001394   0.7703147052576124   0.9801080687388835   0.7568300268401709   0.9001272938154031   0.6301251148774086   0.6199902085264796   0.09833608356466608   0.024387817756960774   0.12237873392320779   0.436727193181721   0.10586600583019369   0.9631256800532806   0.01172968513039126   0.5374708545579379   0.13640647899246883   0.5645357106315863   0.11319118789510511   0.8706958094304192   0.638057065474493   0.3432100499582674   0.9589664700831249   0.08788134242987797   0.3991431054132323   0.5535657116581281   0.1886517648255125   0.10777327369099456   0.6423130785730614   0.6534384178427248   0.5585266499481039   0.48778306516451503   0.5439769950083954   0.6290506000857641   0.4361479160248961   0.051055871982794   0.4381109891782016   0.6659249200324835   0.4244182308945048   0.5135850174248562   0.3017045101857328   0.10138920940089732   0.31122704299939974   0.6428892079944369   0.6636474447112398   0.7581791594426298   0.35226057291627483
0.5550078655645589   0.2645043392980075   0.20461344778450183   0.16360880809076236   0.44723459187356446   0.6221912607249461   0.5511750299417769   0.6050821581426585   0.9594515267090494   0.0782142657165508   0.9221244298560128   0.1689342421177624   0.9083956547262554   0.6401032765383492   0.25619950982352935   0.7445160112232576   0.39481063730139926   0.3383987663526164   0.15481030042263205   0.4332889682238579   0.7519214293069623   0.6747513216413766   0.3966311409800022   0.08102839530758302   0.19691356374240332   0.4102469823433691   0.19201769319550036   0.9174195872168207   0.7496789718688389   0.788055721618423   0.6408426632537234   0.3123374290741622   0.7902274451597894   0.7098414559018722   0.7187182333977105   0.14340318695639978   0.881831790433534   0.06973817936352301   0.46251872357418117   0.3988871757331422   0.48702115313213473   0.7313394130109067   0.3077084231515491   0.9655982075092844   0.7350997238251724   0.05658809136953002   0.9110772821715469   0.8845698122017013   0.5381861600827691   0.6463411090261609   0.7190595889760466   0.9671502249848807   0.7885071882139303   0.8582853874077379   0.0782169257223232   0.6548127959107185   0.9982797430541408   0.14844393150586568   0.3594986923246127   0.5114096089543186   0.11644795262060682   0.07870575214234267   0.8969799687504315   0.11252243322117648
0.6294267994884721   0.34736633913143605   0.5892715455988824   0.14692422571189212   0.8943270756632997   0.29077824776190603   0.6781942634273355   0.2623544135101908   0.35614091558053057   0.6444371387357452   0.9591346744512889   0.29520418852531016   0.5676337273666003   0.7861517513280072   0.8809177487289657   0.6403913926145917   0.5693539843124595   0.6377078198221415   0.521419056404353   0.128981783660273   0.4529060316918527   0.5590020676797989   0.6244390876539215   0.0164593504390965   0.8234792322033806   0.21163572854836282   0.035167542055039074   0.8695351247272044   0.9291521565400809   0.9208574807864568   0.35697327862770356   0.6071807112170136   0.5730112409595502   0.2764203420507117   0.39783860417641465   0.3119765226917034   0.005377513592949973   0.49026859072270446   0.5169208554474489   0.6715851300771117   0.4360235292804905   0.8525607709005629   0.9955017990430959   0.5426033464168387   0.9831174975886378   0.29355870322076405   0.37106271138917446   0.5261439959777423   0.15963826538525722   0.08192297467240123   0.3358951693341354   0.6566088712505379   0.2304861088451763   0.16106549388594443   0.9789218907064318   0.04942816003352433   0.657474867885626   0.8846451518352327   0.5810832865300171   0.737451637341821   0.652097354292676   0.3943765611125283   0.06416243108256815   0.06586650726470918
0.21607382501218558   0.5418157902119654   0.06866063203947223   0.5232631608478704   0.2329563274235478   0.24825708699120125   0.6975979206502978   0.9971191648701282   0.0733180620382906   0.16633411231880002   0.3617027513161624   0.3405102936195903   0.8428319531931142   0.005268618432855601   0.38278086060973066   0.29108213358606594   0.18535708530748823   0.12062346659762287   0.8016975740797135   0.553630496244245   0.5332597310148122   0.7262469054850946   0.7375351429971454   0.4877639889795358   0.31718590600262664   0.18443111527312928   0.6688745109576731   0.9645008281316654   0.08422957857907881   0.9361740282819281   0.9712765903073753   0.9673816632615373   0.010911516540788223   0.769839915963128   0.609573838991213   0.626871369641947   0.16807956334767396   0.7645712975302724   0.2267929783814823   0.33578923605588107   0.9827224780401858   0.6439478309326495   0.4250954043017688   0.7821587398116361   0.44946274702537353   0.9177009254475549   0.6875602613046234   0.2943947508321002   0.1322768410227469   0.7332698101744256   0.01868575034695029   0.32989392270043477   0.048047262443668075   0.7970957818924976   0.04740916003957494   0.3625122594388975   0.03713574590287985   0.0272558659293696   0.43783532104836204   0.7356408897969505   0.8690561825552059   0.2626845683990972   0.2110423426668797   0.3998516537410694
0.8863337045150201   0.6187367374664476   0.785946938365111   0.6176929139294334   0.43687095748964666   0.7010358120188928   0.09838667706048751   0.32329816309733317   0.3045941164668998   0.9677660018444671   0.07970092671353722   0.9934042403968983   0.25654685402323174   0.17067021995196952   0.03229176667396228   0.6308919809580009   0.21941110812035186   0.14341435402259992   0.5944564456256003   0.8952510911610504   0.35035492556514597   0.8807297856235027   0.3834141029587206   0.495399437419981   0.4640212210501258   0.26199304815705504   0.5974671645936096   0.8777065234905476   0.0271502635604791   0.5609572361381623   0.4990804875331221   0.5544083603932145   0.7225561470935793   0.5931912342936952   0.4193795608195849   0.561004119996316   0.46600929307034755   0.4225210143417257   0.3870877941456226   0.9301121390383152   0.2465981849499957   0.27910666031912573   0.7926313485200224   0.03486104787726482   0.8962432593848497   0.39837687469562305   0.4092172455613018   0.5394616104572838   0.43222203833472395   0.13638382653856798   0.8117500809676922   0.6617550869667362   0.40507177477424483   0.5754265904004057   0.31266959343457007   0.1073467265735218   0.6825156276806655   0.9822353561067105   0.8932900326149852   0.5463426065772057   0.21650633461031796   0.5597143417649848   0.5062022384693625   0.6162304675388905
0.9699081496603222   0.28060768144585907   0.7135708899493401   0.5813694196616257   0.07366489027547253   0.882230806750236   0.3043536443880384   0.041907809204341846   0.6414428519407486   0.7458469802116681   0.4926035634203462   0.3801527222376056   0.23637107716650374   0.17042038981126237   0.1799339699857762   0.2728059956640838   0.5538554494858382   0.1881850337045519   0.2866439373707911   0.726463389086878   0.3373491148755203   0.6284706919395671   0.7804416989014286   0.11023292154798754   0.367440965215198   0.34786301049370805   0.06687080895208833   0.5288635018863619   0.29377607493972546   0.46563220374347203   0.7625171645640499   0.48695569268202   0.6523332229989769   0.719785223531804   0.26991360114370366   0.10680297044441439   0.41596214583247315   0.5493648337205417   0.08997963115792747   0.8339969747803306   0.862106696346635   0.36117980001598976   0.8033356937871364   0.10753358569345253   0.5247575814711146   0.7327091080764226   0.022893994885707886   0.997300664145465   0.15731661625591664   0.38484609758271465   0.9560231859336196   0.46843716225910315   0.8635405413161912   0.9192138938392426   0.19350602136956965   0.9814814695770832   0.2112073183172143   0.19942867030743863   0.923592420225866   0.8746784991326687   0.7952451724847411   0.650063836586897   0.8336127890679386   0.040681524352338155
0.9331384761381063   0.2888840365709072   0.030277095280802104   0.9331479386588856   0.4083808946669916   0.5561749284944846   0.007383100395094218   0.9358472745134206   0.251064278411075   0.17132883091176992   0.05135991446147466   0.4674101122543175   0.3875237370948838   0.2521149370725273   0.857853893091905   0.48592864267723435   0.1763164187776695   0.052686266765088675   0.934261472866039   0.6112501435445655   0.3810712462929283   0.40262243017819166   0.10064868379810053   0.5705686191922275   0.447932770154822   0.11373839360728444   0.07037158851729843   0.6374206805333418   0.03955187548783043   0.5575634651127999   0.06298848812220421   0.7015734060199211   0.7884875970767554   0.38623463420102994   0.011628573660729552   0.2341632937656037   0.4009638599818717   0.13411969712850264   0.15377468056882454   0.7482346510883694   0.2246474412042022   0.08143343036341397   0.21951320770278548   0.13698450754380376   0.8435761949112739   0.6788110001852223   0.11886452390468497   0.5664158883515763   0.3956434247564518   0.5650726065779379   0.048492935387386533   0.9289952078182345   0.3560915492686214   0.0075091414651379884   0.9855044472651823   0.22742180179831337   0.5676039521918659   0.621274507264108   0.9738758736044527   0.9932585080327097   0.16664009220999426   0.4871548101356054   0.8201011930356282   0.2450238569443403
0.9419926510057921   0.40572137977219147   0.6005879853328427   0.10803934940053656   0.09841645609451824   0.7269103795869691   0.4817234614281578   0.5416234610489602   0.7027730313380665   0.16183777300903132   0.4332305260407712   0.6126282532307257   0.34668148206944505   0.15432863154389334   0.44772607877558895   0.38520645143241233   0.7790775298775791   0.5330541242797853   0.4738502051711362   0.3919479433997026   0.6124374376675848   0.045899314144179866   0.653749012135508   0.14692408645536234   0.6704447866617927   0.6401779343719884   0.053161026802665184   0.03888473705482577   0.5720283305672745   0.9132675547850192   0.5714375653745074   0.49726127600586556   0.8692552992292081   0.751429781775988   0.13820703933373615   0.8846330227751399   0.522573817159763   0.5971011502320946   0.6904809605581472   0.49942657134272755   0.743496287282184   0.06404702595230932   0.21663075538701107   0.10747862794302489   0.13105884961459913   0.018147711808129456   0.5628817432515031   0.9605545414876625   0.4606140629528064   0.377969777436141   0.509720716448838   0.9216698044328367   0.8885857323855318   0.4647022226511218   0.9382831510743306   0.42440852842697124   0.019330433156323823   0.7132724408751339   0.8000761117405943   0.5397755056518314   0.4967566159965608   0.11617129064303928   0.10959515118244716   0.04034893430910383
0.7532603287143769   0.052124264690729956   0.8929643957954361   0.9328703063660789   0.6222014790997777   0.0339765528826005   0.33008265254393293   0.9723157648784164   0.1615874161469713   0.6560067754464595   0.820361936095095   0.050645960445579605   0.2730016837614394   0.19130455279533765   0.8820787850207644   0.6262374320186084   0.2536712506051156   0.4780321119202038   0.08200267328017007   0.08646192636677699   0.7569146346085548   0.3618608212771645   0.9724075220977229   0.04611299205767316   0.003654305894177981   0.30973655658643456   0.07944312630228681   0.11324268569159422   0.3814528267944003   0.275760003703834   0.7493604737583539   0.14092692081317781   0.21986541064742895   0.6197532282573746   0.9289985376632589   0.09028096036759822   0.9468637268859895   0.4284486754620369   0.046919752642494414   0.4640435283489899   0.6931924762808739   0.9504165635418331   0.9649170793623244   0.37758160198221286   0.9362778416723191   0.5885557422646687   0.9925095572646014   0.3314686099245397   0.9326235357781412   0.2788191856782341   0.9130664309623147   0.21822592423294548   0.5511707089837409   0.0030591819744000713   0.16370595720396078   0.07729900341976766   0.3313052983363119   0.38330595371702547   0.23470741954070193   0.9870180430521694   0.3844415714503224   0.9548572782549886   0.1877876668982075   0.5229745147031796
0.6912490951694484   0.0044407147131554124   0.22287058753588315   0.14539291272096672   0.7549712534971293   0.41588497244848677   0.23036103027128169   0.813924302796427   0.8223477177189882   0.13706578677025266   0.31729459930896703   0.5956983785634815   0.2711770087352473   0.13400660479585258   0.15358864210500625   0.5183993751437138   0.9398717103989354   0.7507006510788271   0.9188812225643044   0.5313813320915445   0.555430138948613   0.7958433728238385   0.7310935556660968   0.008406817388364851   0.8641810437791646   0.7914026581106831   0.5082229681302137   0.8630139046673981   0.10920979028203523   0.37551768566219634   0.277861937858932   0.04908960187097114   0.286862072563047   0.2384518988919437   0.9605673385499649   0.4533912233074896   0.01568506382779971   0.10444529409609112   0.8069786964449587   0.9349918481637758   0.0758133534288643   0.35374464301726405   0.8880974738806543   0.4036105160722313   0.5203832144802513   0.5579012701934255   0.1570039182145575   0.39520369868386646   0.6562021707010868   0.7664986120827424   0.6487809500843438   0.5321897940164684   0.5469923804190515   0.39098092642054605   0.37091901222541185   0.4831001921454972   0.2601303078560045   0.15252902752860234   0.4103516736754469   0.029708968838007582   0.24444524402820478   0.048083733432511204   0.6033729772304882   0.09471712067423183
0.16863189059934044   0.6943390904152472   0.7152755033498339   0.6911066046020005   0.6482486761190892   0.1364378202218217   0.5582715851352764   0.295902905918134   0.9920465054180024   0.36993920813907927   0.9094906350509326   0.7637131119016657   0.4450541249989509   0.9789582817185333   0.5385716228255207   0.2806129197561685   0.18492381714294642   0.826429254189931   0.12821994915007384   0.2509039509181609   0.9404785731147417   0.7783455207574197   0.5248469719195856   0.15618683024392907   0.7718466825154012   0.08400643034217256   0.8095714685697517   0.4650802256419286   0.12359800639631206   0.9475686101203509   0.25129988343447524   0.16917731972379454   0.13155150097830964   0.5776294019812716   0.3418092483835426   0.4054642078221289   0.6864973759793587   0.5986711202627383   0.8032376255580218   0.1248512880659604   0.5015735588364123   0.7722418660728074   0.675017676407948   0.8739473371477995   0.5610949857216706   0.9938963453153876   0.15017070448836242   0.7177605069038704   0.7892483032062694   0.9098899149732151   0.3405992359186108   0.25268028126194186   0.6656502968099574   0.9623213048528643   0.08929935248413555   0.0835029615381473   0.5340987958316477   0.3846919028715926   0.7474901041005929   0.6780387537160184   0.847601419852289   0.7860207826088543   0.9442524785425711   0.553187465650058
0.3460278610158767   0.013778916536046926   0.2692348021346231   0.6792401285022586   0.7849328752942061   0.019882571220659274   0.11906409764626065   0.9614796215983881   0.9956845720879367   0.10999265624744417   0.7784648617276498   0.7087993403364462   0.33003427527797935   0.14767135139457996   0.6891655092435143   0.6252963787982989   0.7959354794463317   0.7629794485229874   0.9416754051429214   0.9472576250822805   0.9483340595940426   0.976958665914133   0.9974229266003503   0.3940701594322225   0.6023061985781659   0.963179749378086   0.7281881244657272   0.714830030929964   0.8173733232839598   0.9432971781574269   0.6091240268194665   0.7533504093315758   0.8216887511960231   0.8333045219099826   0.8306591650918167   0.0445510689951296   0.49165447591804384   0.6856331705154027   0.14149365584830237   0.41925469019683065   0.6957189964717122   0.9226537219924154   0.19981825070538098   0.47199706511455014   0.7473849368776695   0.9456950560782823   0.20239532410503067   0.07792690568232764   0.14507873829950357   0.9825153067001963   0.47420719963930347   0.3630968747523637   0.32770541501554373   0.039218128542769425   0.8650831728198369   0.6097464654207878   0.5060166638195205   0.2059136066327868   0.034424007728020185   0.5651953964256583   0.014362187901476716   0.5202804361173841   0.8929303518797178   0.1459407062288276
0.31864319142976455   0.5976267141249687   0.6931121011743369   0.6739436411142775   0.571258254552095   0.6519316580466864   0.49071677706930616   0.5960167354319498   0.42617951625259143   0.6694163513464901   0.016509577430002708   0.23291986067958612   0.09847410123704772   0.6301982228037207   0.15142640461016582   0.6231733952587982   0.5924574374175272   0.42428461617093394   0.11700239688214564   0.05797799883314002   0.5780952495160505   0.9040041800535499   0.22407204500242783   0.9120372926043124   0.2594520580862859   0.3063774659285811   0.530959943828091   0.23809365149003495   0.6881938035341909   0.6544458078818947   0.04024316675878483   0.6420769160580851   0.2620142872815995   0.9850294565354045   0.023733589328782122   0.40915705537849906   0.16354018604455176   0.3548312337316838   0.8723071847186163   0.7859836601197008   0.5710827486270246   0.9305466175607499   0.7553047878364707   0.7280056612865607   0.9929874991109741   0.026542437507199954   0.5312327428340429   0.8159683686822483   0.7335354410246882   0.7201649715786188   0.0002727990059518315   0.5778747171922134   0.045341637490497265   0.06571916369672416   0.960029632247167   0.9357978011341282   0.7833273502088978   0.08068970716131965   0.9362960429183849   0.5266407457556291   0.619787164164346   0.7258584734296359   0.06398885819976859   0.7406570856359285
0.04870441553732143   0.7953118558688861   0.3086840703632979   0.012651424349367673   0.055716916426347324   0.7687694183616861   0.777451327529255   0.19668305566711936   0.32218147540165915   0.04860444678306728   0.7771785285233033   0.618808338474906   0.2768398379111619   0.9828852830863432   0.8171488962761363   0.6830105373407778   0.4935124877022641   0.9021955759250234   0.8808528533577514   0.15636979158514858   0.8737253235379181   0.17633710249538756   0.8168639951579828   0.41571270594922016   0.8250209080005967   0.3810252466265015   0.5081799247946849   0.4030612815998525   0.7693039915742493   0.6122558282648154   0.7307285972654298   0.20637822593273314   0.4471225161725902   0.5636513814817481   0.9535500687421266   0.5875698874578271   0.17028267826142832   0.5807660983954049   0.13640117246599023   0.9045593501170494   0.6767701905591642   0.6785705224703815   0.25554831910823883   0.7481895585319008   0.8030448670212461   0.5022334199749939   0.438684323950256   0.33247685258268067   0.9780239590206495   0.12120817334849246   0.9305043991555711   0.9294155709828282   0.20871996744640017   0.5089523450836771   0.19977580189014135   0.7230373450500951   0.76159745127381   0.9453009636019291   0.24622573314801485   0.13546745759226794   0.5913147730123817   0.36453486520652406   0.1098245606820246   0.23090810747521853
0.9145445824532175   0.6859643427361426   0.8542762415737858   0.4827185489433177   0.1114997154319713   0.18373092276114864   0.41559191762352976   0.15024169636063703   0.1334757564113218   0.06252274941265616   0.4850875184679586   0.22082612537780882   0.9247557889649216   0.5535704043289791   0.2853117165778173   0.49778878032771373   0.16315833769111168   0.60826944072705   0.03908598342980244   0.3623213227354458   0.57184356467873   0.24373457552052594   0.9292614227477778   0.13141321526022726   0.6572989822255126   0.5577702327843833   0.07498518117399205   0.6486946663169095   0.5457992667935413   0.3740393100232347   0.6593932635504623   0.4984529699562725   0.4123235103822195   0.3115165606105786   0.17430574508250368   0.2776268445784637   0.4875677214172978   0.7579461562815996   0.8889940285046863   0.77983806425075   0.3244093837261861   0.1496767155545495   0.8499080450748839   0.41751674151530416   0.7525658190474561   0.9059421400340235   0.9206466223271061   0.2861035262550769   0.0952668368219435   0.3481719072496402   0.845661441153114   0.6374088599381674   0.5494675700284022   0.9741325972264054   0.18626817760265174   0.13895588998189487   0.13714405964618276   0.6626160366158269   0.011962432520148072   0.8613290454034312   0.6495763382288849   0.9046698803342273   0.12296840401546169   0.08149098115268125
0.3251669545026988   0.7549931647796779   0.27306035894057773   0.6639742396373771   0.5726011354552427   0.8490510247456543   0.35241373661347164   0.3778707133823002   0.4773342986332992   0.5008791174960141   0.5067522954603576   0.7404618534441328   0.9278667286048969   0.5267465202696087   0.32048411785770586   0.601505963462238   0.7907226689587142   0.8641304836537818   0.3085216853375578   0.7401769180588067   0.1411463307298293   0.9594606033195544   0.1855532813220961   0.6586859369061255   0.8159793762271305   0.20446743853987648   0.9124929223815184   0.9947116972687484   0.2433782407718878   0.3554164137942221   0.5600791857680467   0.6168409838864481   0.7660439421385886   0.854537296298208   0.0533268903076891   0.8763791304423154   0.8381772135336917   0.3277907760285993   0.7328427724499832   0.27487316698007747   0.04745454457497742   0.46366029237481754   0.42432108711242544   0.5346962489212707   0.9063082138451481   0.5041996890552631   0.23876780579032936   0.8760103120151452   0.09032883761801763   0.2997322505153867   0.326274883408811   0.8812986147463968   0.8469505968461298   0.9443158367211646   0.7661956976407643   0.26445763085994867   0.08090665470754121   0.08977854042295659   0.7128688073330752   0.38807850041763325   0.24272944117384956   0.7619877643943572   0.9800260348830919   0.11320533343755583
0.19527489659887215   0.29832747201953974   0.5557049477706665   0.5785090845162851   0.288966682753724   0.7941277829642766   0.3169371419803372   0.7024987725011399   0.1986378451357064   0.49439553244888984   0.9906622585715261   0.8212001577547431   0.35168724828957654   0.5500796957277253   0.2244665609307619   0.5567425268947944   0.2707805935820353   0.4603011553047687   0.5115977535976867   0.16866402647716114   0.02805115240818578   0.6983133909104114   0.5315717187145947   0.05545869303960531   0.8327762558093136   0.3999859188908717   0.9758667709439283   0.4769496085233202   0.5438095730555896   0.6058581359265951   0.6589296289635911   0.7744508360221802   0.3451717279198832   0.11146260347770529   0.6682673703920649   0.9532506782674373   0.9934844796303067   0.56138290774998   0.443800809461303   0.3965081513726428   0.7227038860482713   0.10108175244521128   0.9322030558636163   0.22784412489548167   0.6946527336400855   0.40276836153479983   0.40063133714902155   0.17238543185587635   0.8618764778307719   0.0027824426439281456   0.42476456620509334   0.6954358233325562   0.3180669047751823   0.396924306717333   0.7658349372415023   0.9209849873103759   0.972895176855299   0.2854617032396277   0.09756756684943745   0.9677343090429387   0.9794106972249924   0.7240787954896477   0.6537667573881345   0.5712261576702958
0.25670681117672106   0.6229970430444365   0.7215637015245181   0.3433820327748142   0.5620540775366355   0.2202286815096366   0.32093236437549655   0.17099660091893787   0.7001775997058636   0.21744623886570844   0.8961677981704033   0.4755607775863817   0.3821106949306813   0.8205219321483754   0.1303328609289009   0.5545757902760058   0.40921551807538226   0.5350602289087477   0.032765294079463464   0.5868414812330671   0.42980482085038985   0.8109814334191   0.378998536691329   0.015615323562771257   0.17309800967366878   0.18798439037466355   0.6574348351668109   0.672233290787957   0.6110439321370332   0.9677557088650269   0.3365024707913143   0.5012366898690191   0.9108663324311697   0.7503094699993185   0.4403346726209111   0.025675912282637457   0.5287556375004884   0.929787537850943   0.3100018116920102   0.47110012200663165   0.11954011942510614   0.3947273089421953   0.2772365176125467   0.8842586407735645   0.6897352985747163   0.5837458755230953   0.8982379809212178   0.8686433172107932   0.5166372889010475   0.3957614851484318   0.24080314575440684   0.19641002642283623   0.9055933567640142   0.4280057762834048   0.9043006749630925   0.6951733365538171   0.9947270243328445   0.6776963062840863   0.4639660023421815   0.6694974242711796   0.46597138683235617   0.7479087684331432   0.1539641906501713   0.19839730226454796
0.34643126740725   0.3531814594909479   0.8767276730376246   0.31413866149098346   0.6566959688325337   0.7694355839678526   0.9784896921164069   0.4454953442801902   0.1400586799314862   0.37367409881942076   0.737686546362   0.249085317857354   0.23446532316747196   0.945668322536016   0.8333858713989075   0.5539119813035369   0.2397382988346274   0.2679720162519297   0.369419869056726   0.8844145570323574   0.7737669120022712   0.5200632478187864   0.21545567840655472   0.6860172547678094   0.4273356445950212   0.1668817883278385   0.33872800536893016   0.37187859327682593   0.7706396757624875   0.3974462043599859   0.36023831325252326   0.9263832489966357   0.6305809958310012   0.023772105540565136   0.6225517668905233   0.6772979311392817   0.3961156726635293   0.07810378300454916   0.7891658954916158   0.12338594983574483   0.1563773738289019   0.8101317667526196   0.41974602643488973   0.2389713928033875   0.38261046182663067   0.2900685189338331   0.20429034802833504   0.5529541380355781   0.9552748172316095   0.12318673060599461   0.8655623426594049   0.18107554475875218   0.18463514146912194   0.7257405262460087   0.5053240294068816   0.25469229576211644   0.5540541456381206   0.7019684207054435   0.8827722625163584   0.5773943646228347   0.15793847297459132   0.6238646377008944   0.09360636702474265   0.45400841478708986
0.001561099145689406   0.8137328709482748   0.6738603405898529   0.2150370219837024   0.6189506373190587   0.5236643520144417   0.4695699925615179   0.6620828839481243   0.6636758200874493   0.40047762140844717   0.604007649902113   0.4810073391893721   0.47904067861832733   0.6747370951624385   0.09868362049523136   0.22631504342725564   0.9249865329802067   0.9727686744569949   0.21591135797887295   0.648920678804421   0.7670480600056154   0.34890403675610054   0.12230499095413032   0.19491226401733108   0.765486960859926   0.5351711658078256   0.44844465036427744   0.9798752420336287   0.14653632354086724   0.011506813793383912   0.9788746578027595   0.31779235808550443   0.48286050345341797   0.6110291923849368   0.3748670079006466   0.8367850188961323   0.003819824835090595   0.9362920972224983   0.2761833874054152   0.6104699754688767   0.07883329185488389   0.9635234227655034   0.06027202942654225   0.9615492966644558   0.3117852318492685   0.6146193860094028   0.9379670384724119   0.7666370326471247   0.5462982709893425   0.07944822020157716   0.48952238810813453   0.7867617906134959   0.39976194744847526   0.06794140640819324   0.510647730305375   0.46896943252799156   0.9169014439950574   0.4569122140232565   0.1357807224047284   0.6321844136318592   0.9130816191599667   0.5206201168007581   0.8595973349993132   0.0217144381629825
0.8342483273050828   0.5570966940352549   0.7993253055727709   0.06016514149852676   0.5224630954558144   0.9424773080258521   0.861358267100359   0.29352810885140207   0.9761648244664718   0.8630290878242749   0.3718358789922245   0.5067663182379061   0.5764028770179965   0.7950876814160817   0.8611881486868496   0.037796885709914595   0.6595014330229393   0.3381754673928251   0.7254074262821211   0.4056124720780554   0.7464198138629726   0.817555350592067   0.865810091282808   0.3838980339150729   0.9121714865578897   0.2604586565568121   0.06648478571003695   0.3237328924165461   0.3897083911020754   0.3179813485309601   0.20512651860967793   0.030204783565144038   0.4135435666356036   0.45495226070668526   0.8332906396174534   0.5234384653272379   0.837140689617607   0.6598645792906036   0.972102490930604   0.4856415796173233   0.17763925659466773   0.3216891118977785   0.24669506464848281   0.08002910753926791   0.43121944273169516   0.5041337613057115   0.3808849733656749   0.696131073624195   0.5190479561738054   0.24367510474889945   0.314400187655638   0.3723981812076489   0.12933956507173   0.9256937562179394   0.10927366904596003   0.34219339764250484   0.7157959984361264   0.4707414955112541   0.2759830294285066   0.818754932315267   0.8786553088185194   0.8108769162206505   0.3038805384979027   0.3331133526979436
0.7010160522238517   0.48918780432287196   0.057185473849419875   0.2530842451586757   0.2697966094921565   0.9850540430171604   0.676300500483745   0.5569531715344807   0.7507486533183512   0.741378938268261   0.36190031282810703   0.1845549903268318   0.6214090882466211   0.8156851820503216   0.25262664378214694   0.842361592684327   0.9056130898104947   0.34494368653906754   0.9766436143536403   0.023606660369060017   0.02695778099197532   0.534066770318417   0.6727630758557377   0.6904933076711164   0.32594172876812366   0.044878965995545056   0.6155776020063178   0.43740906251244066   0.05614511927596711   0.05982492297838463   0.9392771015225728   0.88045589097796   0.305396465957616   0.31844598471012364   0.5773767886944658   0.6959009006511282   0.6839873777109948   0.502760802659802   0.32475014491231885   0.8535393079668012   0.7783742879005001   0.15781711612073454   0.3481065305586785   0.8299326475977412   0.7514165069085248   0.6237503458023175   0.6753434547029408   0.13943933992662483   0.4254747781404012   0.5788713798067724   0.059765852696623004   0.7020302774141841   0.3693296588644341   0.5190464568283878   0.12048875117405015   0.8215743864362242   0.06393319290681808   0.20060047211826415   0.5431119624795843   0.12567348578509596   0.3799458151958232   0.6978396694584621   0.21836181756726544   0.27213417781829474
0.601571527295323   0.5400225533377275   0.8702552870085869   0.44220153022055353   0.8501550203867982   0.91627220753541   0.19491183230564613   0.3027621902939287   0.4246802422463971   0.33740082772863766   0.1351459796090231   0.6007319128797446   0.05535058338196303   0.8183543709002499   0.014657228434972955   0.7791575264435204   0.991417390475145   0.6177538987819857   0.47154526595538865   0.6534840406584245   0.6114715752793217   0.9199142293235236   0.2531834483881232   0.3813498628401297   0.00990004798399865   0.37989167598579604   0.3829281613795363   0.9391483326195762   0.15974502759720038   0.46361946845038593   0.18801632907389015   0.6363861423256475   0.7350647853508033   0.1262186407217483   0.05287034946486703   0.03565422944590291   0.6797142019688402   0.30786426982149845   0.038213121029894076   0.2564967030023825   0.6882968114936953   0.6901103710395128   0.5666678550745055   0.603012662343958   0.07682523621437355   0.7701961417159892   0.3134844066863822   0.22166279950382836   0.06692518823037491   0.3903044657301931   0.930556245306846   0.2825144668842522   0.9071801606331745   0.9266849972798072   0.7425399162329558   0.6461283245586047   0.17211537528237125   0.8004663565580589   0.6896695667680888   0.6104740951127018   0.492401173313531   0.4926020867365604   0.6514564457381947   0.3539773921103193
0.8041043618198357   0.8024917156970477   0.08478859066368928   0.7509647297663612   0.7272791256054622   0.03229557398105852   0.771304183977307   0.5293019302625329   0.6603539373750872   0.6419911082508654   0.840747938670461   0.2467874633782807   0.7531737767419127   0.7153061109710582   0.09820802243750526   0.600659138819676   0.5810584014595415   0.9148397544129993   0.4085384556694165   0.9901850437069742   0.08865722814601046   0.42223766767643883   0.7570820099312218   0.6362076515966549   0.28455286632617477   0.6197459519793912   0.6722934192675325   0.8852429218302936   0.5572737407207126   0.5874503779983327   0.9009892352902255   0.35594099156776077   0.8969198033456254   0.9454592697474673   0.06024129661976434   0.10915352818948008   0.14374602660371266   0.23015315877640907   0.962033274182259   0.5084943893698041   0.5626876251441713   0.31531340436340977   0.5534948185128427   0.5183093456628299   0.47403039699816074   0.8930757366869709   0.7964128085816209   0.882101694066175   0.18947753067198597   0.2733297847075798   0.12411938931408838   0.9968587722358814   0.6322037899512734   0.6858794067092472   0.22313015402386296   0.6409177806681206   0.735283986605648   0.7404201369617799   0.1628888574040986   0.5317642524786405   0.5915379600019354   0.5102669781853708   0.20085558322183955   0.023269863108836365
0.028850334857764115   0.19495357382196105   0.647360764708997   0.5049605174460065   0.5548199378596034   0.3018778371349901   0.8509479561273761   0.6228588233798314   0.3653424071876174   0.028548052427410292   0.7268285668132877   0.6260000511439501   0.733138617236344   0.34266864571816313   0.5036984127894247   0.9850822704758295   0.997854630630696   0.6022485087563832   0.34080955538532615   0.4533180179971891   0.40631667062876076   0.09198153057101241   0.1399539721634866   0.43004815488835274   0.37746633577099664   0.8970279567490513   0.49259320745448965   0.9250876374423462   0.8226463979113933   0.5951501196140613   0.6416452513271136   0.30222881406251484   0.45730399072377587   0.566602067186651   0.9148166845138258   0.6762287629185647   0.7241653734874318   0.22393342146848785   0.41111827172440113   0.6911464924427352   0.7263107428567358   0.6216849127121046   0.07030871633907497   0.23782847444554606   0.319994072227975   0.5297033821410922   0.9303547441755884   0.8077803195571933   0.9425277364569784   0.6326754253920408   0.43776153672109874   0.8826926821148471   0.11988133854558514   0.037525305777979544   0.7961162853939852   0.5804638680523322   0.6625773478218093   0.47092323859132856   0.8812996008801594   0.9042351051337675   0.9384119743343775   0.24698981712284068   0.4701813291557582   0.21308861269103235
0.21210123147764173   0.625304904410736   0.39987261281668324   0.9752601382454863   0.8921071592496667   0.09560152226964384   0.46951786864109485   0.167479818688293   0.9495794227926884   0.462926096877603   0.03175633191999612   0.28478713657344595   0.8296980842471031   0.4254007910996235   0.23564004652601095   0.7043232685211138   0.16712073642529388   0.9544775525082949   0.3543404456458516   0.8000881633873462   0.2287087620909164   0.7074877353854542   0.8841591164900934   0.5869995506963139   0.016607530613274676   0.08218283097471817   0.48428650367341014   0.6117394124508275   0.12450037136360798   0.9865813087050743   0.014768635032315292   0.44425959376253454   0.17492094857091967   0.5236552118274713   0.9830123031123191   0.1594724571890886   0.3452228643238165   0.09825442072784786   0.7473722565863082   0.4551491886679748   0.17810212789852262   0.14377686821955296   0.39303181094045664   0.6550610252806286   0.9493933658076062   0.4362891328340987   0.5088726944503632   0.06806147458431466   0.9327858351943316   0.3541063018593805   0.024586190776953062   0.4563220621334871   0.8082854638307235   0.3675249931543062   0.00981755574463777   0.012062468370952517   0.6333645152598039   0.8438697813268349   0.0268052526323186   0.852590011181864   0.2881416509359874   0.745615360598987   0.27943299604601035   0.3974408225138891
0.1100395230374648   0.6018384923794341   0.8864011851055538   0.7423797972332605   0.1606461572298586   0.16554935954533537   0.37752849065519056   0.6743183226489459   0.22786032203552703   0.8114430576859548   0.3529422998782375   0.2179962605154588   0.4195748582048035   0.4439180645316486   0.3431247441335997   0.2059337921445063   0.7862103429449996   0.6000482832048137   0.3163194915012811   0.35334378096264235   0.49806869200901216   0.8544329226058267   0.03688649545527074   0.9559029584487533   0.3880291689715474   0.25259443022639255   0.150485310349717   0.2135231612154927   0.2273830117416888   0.08704507068105721   0.7729568196945265   0.5392048385665468   0.9995226897061618   0.2756020129951024   0.42001451981628896   0.321208578051088   0.5799478315013583   0.8316839484634538   0.07688977568268926   0.1152747859065817   0.7937374885563587   0.2316356652586401   0.7605702841814082   0.7619310049439394   0.2956687965473465   0.37720274265281345   0.7236837887261374   0.8060280464951861   0.9076396275757992   0.12460831242642088   0.5731984783764205   0.5925048852796934   0.6802566158341103   0.03756324174536368   0.800241658681894   0.05330004671314659   0.6807339261279487   0.7619612287502613   0.380227138865605   0.7320914686620585   0.1007860946265904   0.9302772802868075   0.30333736318291576   0.6168166827554769
0.3070486060702317   0.6986416150281674   0.5427670790015076   0.8548856778115376   0.011379809522885176   0.3214388723753539   0.8190832902753702   0.048857631316351444   0.10374018194708601   0.19683055994893303   0.24588481189894976   0.45635274603665804   0.4234835661129756   0.15926731820356935   0.4456431532170558   0.40305269932351145   0.742749639985027   0.3973060894533081   0.06541601435145077   0.6709612306614529   0.6419635453584366   0.4670288091665006   0.762078651168535   0.054144547905976   0.33491493928820487   0.7683871941383332   0.2193115721670274   0.19925887009443846   0.3235351297653197   0.44694832176297933   0.4002282818916572   0.150401238778087   0.2197949478182337   0.25011776181404627   0.15434346999270745   0.694048492741429   0.7963113817052581   0.09085044361047695   0.7087003167756517   0.2909957934179175   0.0535617417202311   0.6935443541571689   0.6432843024242009   0.6200345627564646   0.4115981963617945   0.2265155449906683   0.8812056512556659   0.5658900148504886   0.07668325707358967   0.4581283508523351   0.6618940790886385   0.3666311447560502   0.75314812730827   0.011180029089355774   0.2616657971969813   0.21622990597796315   0.5333531794900364   0.7610622672753095   0.10732232720427383   0.5221814132365342   0.7370417977847783   0.6702118236648326   0.39862201042862216   0.23118561981861668
0.6834800560645471   0.9766674695076637   0.7553377080044212   0.6111510570621521   0.2718818597027526   0.7501519245169953   0.8741320567487554   0.04526104221166343   0.19519860262916294   0.29202357366466025   0.21223797766011687   0.6786298974556133   0.4420504753208929   0.28084354457530447   0.9505721804631356   0.4623999914776501   0.9086972958308567   0.519781277299995   0.8432498532588618   0.9402185782411159   0.1716554980460784   0.8495694536351625   0.44462784283023965   0.7090329584224992   0.48817544198153123   0.8729019841274989   0.6892901348258184   0.09788190136034713   0.21629358227877865   0.12275005961050348   0.815158078077063   0.0526208591486837   0.021094979649615726   0.8307264859458432   0.6029201004169461   0.37399096169307045   0.5790445043287228   0.5498829413705387   0.6523479199538105   0.9115909702154203   0.6703472084978661   0.030101664070543755   0.8090980666949488   0.9713723919743045   0.49869171045178773   0.18053221043538129   0.36447022386470906   0.2623394335518053   0.01051626847025648   0.30763022630788245   0.6751800890388907   0.16445753219145812   0.7942226861914778   0.184880166697379   0.8600220109618277   0.1118366730427744   0.7731277065418621   0.35415368075153575   0.25710191054488163   0.737845711349704   0.19408320221313932   0.804270739380997   0.6047539905910712   0.8262547411342837
0.5237359937152731   0.7741690753104533   0.7956559238961224   0.8548823491599792   0.025044283263485442   0.593636864875072   0.4311857000314133   0.5925429156081738   0.014528014793228962   0.2860066385671895   0.7560056109925226   0.42808538341671576   0.22030532860175114   0.1011264718698105   0.8959836000306949   0.31624871037394137   0.44717762205988904   0.7469727911182747   0.6388816894858133   0.5784029990242374   0.25309441984674974   0.9427020517372777   0.03412769889474211   0.7521482578899538   0.7293584261314765   0.16853297642682444   0.23847177499861968   0.8972659087299747   0.7043141428679911   0.5748961115517525   0.8072860749672064   0.3047229931218008   0.6897861280747621   0.28888947298456297   0.05128046397468378   0.876637609705085   0.46948079947301097   0.18776300111475247   0.15529686394398892   0.5603888993311437   0.022303177413121954   0.4407902099964777   0.5164151744581756   0.9819859003069062   0.7692087575663722   0.49808815825920005   0.4822874755634336   0.2298376424169524   0.0398503314348957   0.3295551818323756   0.2438157005648139   0.33257173368697773   0.3355361885669046   0.7546590702806231   0.4365296255976075   0.02784874056517696   0.6457500604921425   0.46576959729606016   0.3852491616229237   0.15121113086009197   0.17626926101913148   0.2780065961813077   0.2299522976789348   0.5908222315289483
0.15396608360600952   0.83721638618483   0.7135371232207591   0.6088363312220422   0.3847573260396373   0.3391282279256299   0.23124964765732553   0.37899868880508975   0.3449069946047416   0.00957304609325433   0.9874339470925116   0.04642695511811204   0.00937080603783699   0.2549139758126312   0.5509043214949041   0.01857821455293508   0.3636207455456945   0.789144378516571   0.16565515987198043   0.8673670836928431   0.18735148452656303   0.5111377823352634   0.9357028621930457   0.27654485216389474   0.0333854009205535   0.6739213961504334   0.2221657389722865   0.6677085209418526   0.6486280748809162   0.33479316822480354   0.990916091314961   0.2887098321367628   0.3037210802761746   0.3252201221315492   0.003482144222449338   0.24228287701865078   0.2943502742383376   0.07030614631891799   0.4525778227275452   0.22370466246571571   0.9307295286926431   0.2811617678023469   0.2869226628555648   0.3563375787728726   0.7433780441660801   0.7700239854670835   0.3512198006625191   0.07979272660897785   0.7099926432455266   0.0961025893166501   0.12905406169023262   0.4120842056671253   0.06136456836461038   0.7613094210918466   0.13813797037527165   0.12337437353036244   0.7576434880884357   0.43608929896029736   0.13465582615282232   0.8810914965117117   0.46329321385009814   0.3657831526413794   0.6820780034252771   0.657386834045996
0.5325636851574551   0.08462138483903248   0.39515534056971235   0.3010492552731234   0.789185640991375   0.3145973993719489   0.04393553990719319   0.22125652866414552   0.07919299774584841   0.21849481005529883   0.9148814782169605   0.8091723229970202   0.017828429381238037   0.4571853889634523   0.7767435078416889   0.6857979494666578   0.2601849412928023   0.02109609000315489   0.6420876816888667   0.8047064529549461   0.7968917274427041   0.6553129373617755   0.9600096782635895   0.1473196189089502   0.26432804228524903   0.5706915525227431   0.5648543376938772   0.8462703636358269   0.47514240129387403   0.2560941531507941   0.5209187977866839   0.6250138349716813   0.39594940354802566   0.03759934309549523   0.6060373195697234   0.815841511974661   0.3781209741667876   0.580413954132043   0.8292938117280345   0.13004356250800325   0.11793603287398532   0.5593178641288881   0.18720613003916786   0.3253371095530571   0.3210443054312812   0.9040049267671125   0.22719645177557837   0.17801749064410688   0.05671626314603219   0.3333133742443696   0.6623421140817012   0.3317471270082801   0.5815738618521581   0.07721922109357549   0.14142331629501723   0.7067332920365987   0.18562445830413252   0.039619877998080255   0.5353859967252939   0.8908917800619377   0.807503484137345   0.4592059238660373   0.7060921849972593   0.7608482175539344
0.6895674512633596   0.8998880597371492   0.5188860549580915   0.43551110800087733   0.36852314583207835   0.9958831329700366   0.2916896031825131   0.2574936173567704   0.31180688268604617   0.6625697587256671   0.6293474891008118   0.9257464903484903   0.7302330208338881   0.5853505376320917   0.4879241728057947   0.21901319831189164   0.5446085625297555   0.5457306596340114   0.9525381760805008   0.328121418249954   0.7371050783924106   0.08652473576797406   0.24644599108324156   0.5672732006960196   0.04753762712905104   0.18663667603082484   0.7275599361251501   0.13176209269514225   0.6790144812969727   0.19075354306078818   0.43587033294263705   0.8742684753383718   0.3672075986109265   0.528183784335121   0.8065228438418252   0.9485219849898815   0.6369745777770385   0.9428332467030295   0.3185986710360305   0.7295087866779898   0.09236601524728297   0.39710258706901813   0.3660604949555296   0.40138736842803585   0.35526093685487237   0.31057785130104404   0.11961450387228806   0.8341141677320163   0.3077233097258213   0.12394117527021922   0.3920545677471379   0.702352075036874   0.6287088284288487   0.933187632209431   0.9561842348045009   0.8280835996985022   0.2615012298179221   0.40500384787430993   0.14966139096267572   0.8795616147086208   0.6245266520408836   0.4621706011712805   0.8310627199266453   0.15005282803063094
0.5321606367936007   0.06506801410226236   0.46500222497111565   0.7486654596025951   0.1768996999387283   0.7544901628012183   0.3453877210988276   0.9145512918705788   0.869176390212907   0.6305489875309991   0.9533331533516897   0.21219921683370482   0.24046756178405837   0.6973613553215681   0.9971489185471888   0.3841156171352026   0.9789663319661362   0.2923575074472581   0.8474875275845131   0.5045540024265819   0.35443967992525266   0.8301869062759776   0.016424807657867767   0.35450117439595086   0.822279043131652   0.7651188921737152   0.5514225826867521   0.6058357147933557   0.6453793431929237   0.010628729372496938   0.20603486158792456   0.6912844229227769   0.7762029529800167   0.38007974184149784   0.2527017082362349   0.4790852060890721   0.5357353911959584   0.6827183865199298   0.25555278968904616   0.0949695889538695   0.556769059229822   0.3903608790726717   0.40806526210453314   0.5904155865272877   0.2023293793045694   0.5601739727966941   0.39164045444666534   0.2359144121313368   0.3800503361729174   0.7950550806229789   0.8402178717599132   0.630078697337981   0.7346709929799937   0.7844263512504819   0.6341830101719886   0.9387942744152041   0.958468039999977   0.4043466094089841   0.3814813019357538   0.459709068326132   0.4227326488040187   0.7216282228890543   0.12592851224670762   0.36473947937226253
0.8659635895741966   0.33126734381638256   0.7178632501421744   0.7743238928449748   0.6636342102696272   0.7710933710196884   0.3262227956955091   0.538409480713638   0.2835838740967098   0.9760382903967095   0.4860049239355959   0.908330783375657   0.5489128811167162   0.19161193914622765   0.8518219137636072   0.9695365089604528   0.5904448411167391   0.7872653297372436   0.4703406118278534   0.5098274406343208   0.1677121923127205   0.06563710684818931   0.3444120995811458   0.1450879612620583   0.3017486027385239   0.7343697630318068   0.6265488494389713   0.3707640684170835   0.6381143924688967   0.9632763920121183   0.3003260537434622   0.8323545877034454   0.3545305183721868   0.9872381016154087   0.8143211298078663   0.9240238043277884   0.8056176372554706   0.7956261624691812   0.9624992160442591   0.9544872953673356   0.21517279613873147   0.008360832731937533   0.49215860421640567   0.4446598547330147   0.04746060382601097   0.9427237258837482   0.14774650463525987   0.2995718934709564   0.7457120010874871   0.20835396285194147   0.5211976551962886   0.9288078250538729   0.10759760861859044   0.24507757083982312   0.22087160145282636   0.09645323735042749   0.7530670902464036   0.25783946922441436   0.40655047164496005   0.17242943302263905   0.947449452990933   0.46221330675523326   0.44405125560070097   0.2179421376553035
0.7322766568522016   0.4538524740232957   0.9518926513842952   0.7732822829222887   0.6848160530261905   0.5111287481395475   0.8041461467490354   0.47371038945133237   0.9391040519387035   0.30277478528760604   0.2829484915527468   0.5449025643974594   0.831506443320113   0.05769721444778292   0.06207689009992045   0.44844932704703194   0.07843935307370939   0.7998577452233685   0.6555264184549604   0.27601989402439286   0.1309899000827764   0.3376444384681353   0.21147516285425944   0.058077756369089385   0.3987132432305749   0.8837919644448395   0.25958251146996414   0.2847954734468006   0.7138971902043844   0.37266321630529203   0.4554363647209288   0.8110850839954683   0.7747931382656809   0.069888431017686   0.17248787316818195   0.2661825195980088   0.9432866949455679   0.012191216569903088   0.1104109830682615   0.8177331925509769   0.8648473418718585   0.21233347134653455   0.4548845646133011   0.541713298526584   0.7338574417890821   0.8746890328783993   0.2434094017590417   0.4836355421574946   0.3351441985585072   0.9908970684335597   0.9838268902890775   0.198840068710694   0.6212470083541228   0.6182338521282676   0.5283905255681487   0.38775498471522574   0.846453870088442   0.5483454211105816   0.35590265239996677   0.12157246511721691   0.903167175142874   0.5361542045406785   0.2454916693317053   0.30383927256624
0.038319833271015555   0.323820733194144   0.7906071047184042   0.762125974039656   0.30446239148193344   0.44913170031574473   0.5471977029593625   0.2784904318821614   0.9693181929234262   0.45823463188218505   0.563370812670285   0.07965036317146736   0.3480711845693034   0.8400007797539174   0.03498028710213626   0.6918953784562416   0.5016173144808614   0.2916553586433358   0.6790776347021694   0.5703229133390247   0.5984501393379874   0.7555011541026573   0.4335859653704642   0.2664836407727847   0.5601303060669719   0.4316804209085133   0.64297886065206   0.5043576667331287   0.2556679145850384   0.9825487205927685   0.0957811576926975   0.22586723485096732   0.28634972166161216   0.5243140887105835   0.5324103450224125   0.14621687167949998   0.9382785370923088   0.6843133089566661   0.4974300579202763   0.4543214932232584   0.4366612226114473   0.39265795031333023   0.8183524232181068   0.8839985798842337   0.83821108327346   0.637156796210673   0.38476645784764263   0.617514939111449   0.27808077720648805   0.2054763753021597   0.7417875971955826   0.11315727237832025   0.022412862621449665   0.2229276547093912   0.646006439502885   0.8872900375273529   0.7360631409598375   0.6986135659988078   0.11359609448047259   0.741073165847853   0.7977846038675288   0.014300257042141695   0.6161660365601963   0.28675167262459456
0.3611233812560815   0.6216423067288115   0.7978136133420896   0.4027530927403609   0.5229122979826216   0.9844855105181385   0.4130471554944469   0.785238153628912   0.24483152077613354   0.7790091352159788   0.6712595582988643   0.6720808812505917   0.22241865815468387   0.5560814805065876   0.02525311879597925   0.7847908437232388   0.4863555171948464   0.8574679145077798   0.9116570243155067   0.04371767787538586   0.6885709133273176   0.8431676574656382   0.29549098775531035   0.7569660052507913   0.3274475320712361   0.22152535073682672   0.4976773744132208   0.35421291251043036   0.8045352340886145   0.2370398402186882   0.08463021891877384   0.5689747588815184   0.5597037133124809   0.4580307050027094   0.4133706606199095   0.8968938776309267   0.3372850551577971   0.9019492244961218   0.38811754182393027   0.11210303390768785   0.8509295379629508   0.044481309988341974   0.4764605175084236   0.06838535603230199   0.16235862463563316   0.2013136525227038   0.18096952975311326   0.31141935078151073   0.8349110925643971   0.9797883017858771   0.6832921553398924   0.9572064382710803   0.03037585847578258   0.7427484615671889   0.5986619364211186   0.388231679389562   0.47067214516330164   0.28471775656447945   0.1852912758012091   0.49133780175863534   0.13338709000550453   0.3827685320683576   0.7971737339772789   0.3792347678509475
0.28245755204255374   0.33828722208001566   0.32071321646885526   0.3108494118186455   0.12009892740692059   0.13697356955731183   0.13974368671574203   0.9994300610371348   0.2851878348425235   0.15718526777143474   0.45645153137584954   0.042223622766054444   0.2548119763667409   0.41443680620424583   0.857789594954731   0.6539919433764925   0.7841398312034393   0.1297190496397664   0.6724983191535219   0.16265414161785707   0.6507527411979348   0.7469505175714088   0.875324585176243   0.7834193737669096   0.36829518915538106   0.4086632954913932   0.5546113687073877   0.47256996194826406   0.24819626174846043   0.27168972593408136   0.4148676819916457   0.47313990091112923   0.9630084269059369   0.11450445816264661   0.9584161506157961   0.43091627814507477   0.708196450539196   0.7000676519584007   0.1006265556610652   0.7769243347685824   0.9240566193357567   0.5703486023186344   0.42812823650754334   0.6142701931507253   0.27330387813782187   0.8233980847472255   0.5528036513313004   0.8308508193838157   0.9050086889824408   0.4147347892558324   0.9981922826239127   0.35828085743555166   0.6568124272339804   0.14304506332175107   0.583324600632267   0.8851409565244224   0.6938040003280435   0.028540605159104462   0.6249084500164708   0.45422467837934766   0.9856075497888475   0.3284729532007037   0.5242818943554056   0.6773003436107653
0.06155093045309076   0.7581243508820693   0.09615365784786226   0.06303015046004001   0.7882470523152689   0.9347262661348438   0.5433500065165618   0.23217933107622432   0.883238363332828   0.5199914768790114   0.5451577238926493   0.8738984736406726   0.22642593609884765   0.37694641355726033   0.9618331232603823   0.9887575171162503   0.5326219357708042   0.3484058083981558   0.3369246732439115   0.5345328387369026   0.5470143859819567   0.019932855197452144   0.8126427788885059   0.8572324951261373   0.48546345552886594   0.2618085043153828   0.7164891210406437   0.7942023446660973   0.6972164032135971   0.327082238180539   0.17313911452408176   0.5620230135898729   0.813978039880769   0.8070907613015277   0.6279813906314325   0.6881245399492003   0.5875521037819214   0.4301443477442673   0.6661482673710502   0.69936702283295   0.054930168011117234   0.08173853934611147   0.3292235941271387   0.1648341840960475   0.5079157820291605   0.06180568414865932   0.5165808152386328   0.3076016889699102   0.022452326500294557   0.7999971798332766   0.8000916941979891   0.5133993443038128   0.3252359232866975   0.4729149416527375   0.6269525796739074   0.9513763307139399   0.5112578834059285   0.6658241803512098   0.9989711890424748   0.26325179076473953   0.923705779624007   0.23567983260694256   0.3328229216714247   0.5638847679317894
0.8687756116128899   0.15394129326083109   0.0035993275442860176   0.39905058383574193   0.3608598295837293   0.09213560911217178   0.48701851230565324   0.09144889486583178   0.33840750308343476   0.2921384292788953   0.6869268181076641   0.5780495505620189   0.013171579796737257   0.8192234876261577   0.05997423843375671   0.626673219848079   0.5019136963908089   0.15339930727494788   0.06100304939128182   0.3634214290833395   0.5782079167668017   0.9177194746680053   0.7281801277198571   0.7995366611515501   0.709432305153912   0.7637781814071742   0.7245808001755711   0.4004860773158081   0.34857247557018267   0.6716425722950025   0.23756228786991787   0.3090371824499763   0.010164972486747937   0.3795041430161072   0.5506354697622537   0.7309876318879575   0.9969933926900106   0.5602806553899494   0.49066123132849704   0.10431441203987837   0.49507969629920184   0.40688134811500154   0.4296581819372152   0.7408929829565388   0.9168717795324001   0.48916187344699624   0.7014780542173581   0.9413563218049888   0.20743947437848811   0.725383692039822   0.976897254041787   0.5408702444891808   0.8588669988083054   0.053741119744819606   0.7393349661718691   0.2318330620392044   0.8487020263215576   0.6742369767287124   0.18869949640961536   0.5008454301512469   0.8517086336315468   0.11395632133876302   0.6980382650811183   0.3965310181113686
0.35662893733234496   0.7070749732237614   0.26838008314390305   0.6556380351548298   0.43975715779994484   0.2179130997767652   0.566902028926545   0.7142817133498409   0.23231768342145676   0.4925294077369432   0.590004774884758   0.1734114688606602   0.3734506846131513   0.43878828799212355   0.8506698087128889   0.9415784068214558   0.5247486582915938   0.7645513112634111   0.6619703123032735   0.44073297667020883   0.673040024660047   0.6505949899246481   0.9639320472221552   0.0442019585588402   0.316411087327702   0.9435200167008867   0.6955519640782521   0.38856392340401047   0.8766539295277571   0.7256069169241215   0.12864993515170717   0.6742822100541696   0.6443362461063004   0.23307750918717826   0.5386451602669492   0.5008707411935094   0.2708855614931491   0.7942892211950547   0.6879753515540603   0.5592923343720536   0.7461369032015552   0.029737909931643554   0.026005039250786857   0.11855935770184477   0.07309687854150831   0.37914292000699545   0.06207299202863167   0.07435739914300456   0.7566857912138063   0.43562290330610876   0.36652102795037955   0.6857934757389941   0.8800318616860492   0.7100159863819874   0.23787109279867238   0.011511265684824525   0.23569561557974875   0.4769384771948091   0.6992259325317232   0.5106405244913151   0.9648100540865996   0.6826492559997543   0.011250580977662857   0.9513481901192615
0.21867315088504435   0.6529113460681109   0.985245541726876   0.8327888324174169   0.14557627234353604   0.2737684260611154   0.9231725496982444   0.7584314332744122   0.38889048112972974   0.8381455227550066   0.5566515217478648   0.07263795753541816   0.5088586194436806   0.12812953637301927   0.3187804289491924   0.06112669185059363   0.2731630038639319   0.6511910591782102   0.6195544964174692   0.5504861673592785   0.30835294977733224   0.9685418031784558   0.6083039154398063   0.5991379772400169   0.08967979889228789   0.315630457110345   0.6230583737129304   0.7663491448226001   0.9441035265487518   0.04186203104922958   0.699885824014686   0.007917711548187859   0.555213045419022   0.20371650829422297   0.1432343022668212   0.9352797540127697   0.04635442597534148   0.07558697192120367   0.8244538733176289   0.874153062162176   0.7731914221114096   0.4243959127429935   0.20489937690015966   0.3236668948028976   0.4648384723340774   0.45585410956453765   0.5965954614603534   0.7245289175628807   0.3751586734417895   0.14022365245419266   0.973537087747423   0.9581797727402805   0.43105514689303764   0.09836162140496309   0.273651263732737   0.9502620611920928   0.8758421014740155   0.8946451131107401   0.13041696146591578   0.014982307179323029   0.8294876754986741   0.8190581411895365   0.30596308814828693   0.14082924501714694
0.05629625338726448   0.394662228446543   0.10106371124812728   0.8171623502142493   0.5914577810531871   0.9388081188820053   0.5044682497877739   0.09263343265136866   0.21629910761139762   0.7985844664278127   0.530931162040351   0.13445365991108804   0.78524396071836   0.7002228450228496   0.257279898307614   0.18419159871899532   0.9094018592443445   0.8055777319121095   0.12686293684169822   0.1692092915396723   0.07991418374567034   0.986519590722573   0.8208998486934113   0.02838004652252534   0.023617930358405863   0.59185736227603   0.719836137445284   0.211217696308276   0.43216014930521873   0.6530492433940246   0.21536788765751003   0.11858426365690734   0.21586104169382112   0.8544647769662119   0.6844367256171591   0.9841306037458193   0.43061708097546114   0.1542419319433624   0.4271568273095451   0.799939005026824   0.5212152217311167   0.3486642000312529   0.3002938904678469   0.6307297134871517   0.44130103798544634   0.36214460930868   0.4793940417744356   0.6023496669646263   0.4176831076270405   0.77028724703265   0.7595579043291516   0.39113197065635036   0.9855229583218218   0.11723800363862531   0.5441900166716416   0.272547706999443   0.7696619166280007   0.2627732266724133   0.8597532910544825   0.2884171032536237   0.3390448356525395   0.10853129472905096   0.43259646374493743   0.4884780982267997
0.8178296139214228   0.759867094697798   0.13230257327709052   0.8577483847396481   0.37652857593597644   0.39772248538911803   0.6529085315026549   0.2553987177750217   0.9588454683089359   0.6274352383564681   0.8933506271735033   0.8642667471186714   0.9733225099871142   0.5101972347178427   0.34916061050186176   0.5917190401192284   0.20366059335911355   0.2474240080454294   0.48940731944737925   0.3033019368656047   0.8646157577065741   0.13889271331637848   0.05681085570244185   0.8148238386388049   0.04678614378515125   0.3790256186185805   0.9245082824253513   0.9570754538991569   0.6702575678491748   0.9813031332294624   0.2715997509226964   0.7016767361241352   0.7114120995402389   0.3538678948729943   0.37824912374919306   0.8374099890054638   0.7380895895531246   0.8436706601551516   0.029088513247331305   0.24569094888623538   0.5344289961940112   0.5962466521097222   0.539681193799952   0.9423890120206307   0.6698132384874371   0.45735393879334363   0.4828703380975102   0.12756517338182577   0.6230270947022858   0.0783283201747632   0.5583620556721589   0.17048971948266886   0.952769526853111   0.09702518694530078   0.28676230474946246   0.4688129833585337   0.24135742731287216   0.7431572920723065   0.9085131810002695   0.6314029943530699   0.5032678377597475   0.8994866319171549   0.8794246677529381   0.3857120454668345
0.9688388415657363   0.3032399798074328   0.3397434739529861   0.44332303344620383   0.29902560307829923   0.8458860410140892   0.8568731358554759   0.31575786006437806   0.6759985083760134   0.7675577208393259   0.298511080183317   0.1452681405817092   0.7232289815229024   0.6705325338940251   0.01174877543385453   0.6764551572231755   0.4818715542100302   0.9273752418217187   0.10323559443358511   0.04505216287010555   0.9786037164502828   0.02788860990456378   0.223810926680647   0.659340117403271   0.00976487488454644   0.724648630097131   0.884067452727661   0.21601708395706717   0.7107392718062472   0.8787625890830418   0.027194316872185046   0.9002592238926891   0.03474076343023387   0.11120486824371591   0.728683236688868   0.75499108331098   0.31151178190733153   0.4406723343496907   0.7169344612550135   0.07853592608780444   0.8296402276973014   0.5132970925279721   0.6136988668214284   0.03348376321769888   0.8510365112470186   0.48540848262340824   0.3898879401407814   0.3741436458144279   0.8412716363624722   0.7607598525262773   0.5058204874131205   0.15812656185736068   0.1305323645562249   0.8819972634432355   0.4786261705409354   0.2578673379646716   0.09579160112599105   0.7707923951995195   0.7499429338520673   0.5028762546536917   0.7842798192186595   0.33012006084982876   0.033008472597053876   0.4243403285658872
0.9546395915213581   0.8168229683218567   0.4193096057756255   0.39085656534818836   0.10360308027433959   0.33141448569844845   0.029421665634844094   0.016712919533760473   0.2623314439118674   0.5706546331721711   0.5236011782217236   0.8585863576763998   0.1317990793556425   0.6886573697289358   0.044975007680788215   0.6007190197117283   0.03600747822965145   0.9178649745294162   0.2950320738287208   0.09784276505803656   0.2517276590109919   0.5877449136795875   0.26202360123166696   0.6735024364921494   0.29708806748963373   0.7709219453577307   0.8427139954560414   0.282645871143961   0.19348498721529414   0.4395074596592823   0.8132923298211974   0.26593295161020053   0.9311535433034267   0.868852826487111   0.28969115159947373   0.40734659393380074   0.7993544639477842   0.18019545675817533   0.24471614391868554   0.8066275742220725   0.7633469857181328   0.2623304822287591   0.9496840700899647   0.708784809164036   0.5116193267071408   0.6745855685491716   0.6876604688582978   0.035282372671886615   0.2145312592175071   0.903663623191441   0.8449464734022563   0.7526365015279256   0.021046272002212933   0.4641561635321587   0.03165414358105891   0.4867035499177251   0.08989272869878621   0.5953033370450476   0.7419629919815852   0.07935695598392434   0.29053826475100203   0.4151078802868723   0.49724684806289965   0.2727293817618518
0.5271912790328692   0.15277739805811316   0.547562777972935   0.5639445725978158   0.015571952325728422   0.4781918295089415   0.8599023091146372   0.5286621999259292   0.8010406931082213   0.5745282063175006   0.014955835712380908   0.7760256983980036   0.7799944211060084   0.11037204278534182   0.983301692131322   0.28932214848027854   0.6901016924072222   0.5150687057402942   0.24133870014973682   0.2099651924963542   0.39956342765622016   0.09996082545342193   0.7440918520868371   0.9372358107345024   0.8723721486233509   0.9471834273953088   0.19652907411390225   0.3732912381366865   0.8568001962976225   0.4689915978863673   0.336626764999265   0.8446290382107573   0.05575950318940118   0.8944633915688668   0.3216709292868841   0.06860333981275368   0.2757650820833928   0.7840913487835249   0.33836923715556216   0.7792811913324751   0.5856633896761706   0.2690226430432307   0.09703053700582531   0.5693159988361209   0.1860999620199504   0.1690618175898088   0.3529386849189881   0.6320801881016186   0.3137278133965995   0.22187839019450004   0.1564096108050859   0.258788949964932   0.45692761709897695   0.7528867923081327   0.8197828458058208   0.4141599117541747   0.4011681139095758   0.858423400739266   0.4981119165189367   0.34555657194142103   0.125403031826183   0.07433205195574107   0.15974267936337455   0.5662753806089459
0.5397396421500125   0.8053094089125103   0.06271214235754922   0.996959381772825   0.35363968013006203   0.6362475913227016   0.7097734574385611   0.3648791936712064   0.03991186673346255   0.4143692011282015   0.5533638466334753   0.10609024370627439   0.5829842496344856   0.6614824088200688   0.7335810008276543   0.6919303319520996   0.1818161357249098   0.8030590080808028   0.23546908430871769   0.34637376001067866   0.05641310389872678   0.7287269561250618   0.07572640494534312   0.7800983794017328   0.5166734617487143   0.9234175472125514   0.013014262587793896   0.7831389976289078   0.1630337816186523   0.28716995588984984   0.3032408051492328   0.41825980395770146   0.12312191488518977   0.8728007547616483   0.7498769585157576   0.31216956025142706   0.5401376652507042   0.21131834594157947   0.016295957688103213   0.6202392282993274   0.3583215295257944   0.40825933786077667   0.7808268733793855   0.2738654682886487   0.3019084256270676   0.679532381735715   0.7051004684340424   0.49376708888691595   0.7852349638783532   0.7561148345231635   0.6920862058462485   0.7106280912580081   0.6222011822597009   0.46894487863331374   0.38884540069701573   0.2923682873003067   0.4990792673745112   0.5961441238716655   0.6389684421812581   0.9801987270488796   0.958941602123807   0.384825777930086   0.6226724844931549   0.3599594987495522
0.6006200725980126   0.9765664400693094   0.8418456111137694   0.08609403046090346   0.298711646970945   0.2970340583335944   0.13674514267972696   0.5923269415739875   0.5134766830925918   0.5409192238104309   0.44465893683347846   0.8816988503159794   0.8912755008328908   0.07197434517711712   0.055813536136462734   0.5893305630156728   0.3921962334583796   0.47583022130545166   0.4168450939552046   0.6091318359667932   0.43325463133457265   0.09100444337536566   0.7941726094620497   0.24917233721724097   0.83263455873656   0.11443800330605633   0.9523269983482803   0.16307830675633753   0.533922911765615   0.8174039449724619   0.8155818556685533   0.57075136518235   0.020446228673023287   0.2764847211620311   0.3709229188350749   0.6890525148663706   0.12917072784013248   0.20451037598491398   0.31510938269861216   0.09972195185069785   0.7369744943817529   0.7286801546794623   0.8982642887434076   0.49059011588390466   0.3037198630471802   0.6376757113040966   0.10409167928135786   0.2414177786666637   0.4710853043106202   0.5232377079980404   0.15176468093307754   0.07833947191032617   0.9371623925450051   0.7058337630255784   0.3361828252645242   0.5075881067279762   0.9167161638719818   0.4293490418635473   0.9652599064294494   0.8185355918616055   0.7875454360318493   0.22483866587863333   0.6501505237308371   0.7188136400109078
0.05057094165009651   0.496158511199171   0.7518862349874297   0.22822352412700306   0.7468510786029163   0.8584827998950744   0.6477945557060718   0.9868057454603394   0.27576577429229615   0.335245091897034   0.4960298747729942   0.9084662735500132   0.33860338174729104   0.6294113288714557   0.15984704950847   0.40087816682203703   0.4218872178753092   0.20006228700790835   0.19458714307902067   0.5823425749604314   0.6343417818434598   0.9752236211292751   0.5444366193481834   0.8635289349495238   0.5837708401933633   0.47906510993010404   0.7925503843607539   0.6353054108225207   0.836919761590447   0.6205823100350297   0.1447558286546821   0.6484996653621813   0.5611539872981508   0.2853372181379957   0.6487259538816879   0.7400333918121681   0.22255060555085981   0.65592588926654   0.4888789043732179   0.3391552249901311   0.8006633876755507   0.4558636022586317   0.2942917612941972   0.7568126500296997   0.1663216058320908   0.48063998112935663   0.7498551419460138   0.8932837150801759   0.5825507656387274   0.0015748711992526333   0.9573047575852599   0.2579783042576553   0.7456310040482804   0.380992561164223   0.8125489289305778   0.6094786388954739   0.18447701675012962   0.09565534302622729   0.1638229750488899   0.8694452470833058   0.9619264111992698   0.43972945375968725   0.674944070675672   0.5302900220931747
0.16126302352371918   0.9838658515010555   0.3806523093814748   0.773477372063475   0.9949414176916284   0.503225870371699   0.6307971674354611   0.8801936569832991   0.41239065205290093   0.5016509991724463   0.6734924098502012   0.6222153527256438   0.6667596480046205   0.12065843800822335   0.8609434809196234   0.012736713830169836   0.48228263125449083   0.025003094981996054   0.6971205058707335   0.14329146674686402   0.5203562200552211   0.5852736412223087   0.02217643519506147   0.6130014446536893   0.3590931965315019   0.6014077897212532   0.6415241258135866   0.8395240725902143   0.3641517788398735   0.09818191934955427   0.010726958378125626   0.9593304156069152   0.9517611267869726   0.596530920177108   0.33723454852792445   0.33711506288127147   0.2850014787823521   0.4758724821688846   0.47629106760830103   0.32437834905110163   0.8027188475278613   0.45086938718688857   0.7791705617375676   0.1810868823042376   0.2823626274726402   0.8655957459645798   0.7569941265425061   0.5680854376505483   0.9232694309411383   0.2641879562433266   0.11547000072891941   0.728561365060334   0.5591176521012649   0.16600603689377233   0.10474304235079379   0.7692309494534187   0.6073565253142923   0.5694751167166644   0.7675084938228693   0.4321158865721472   0.32235504653194014   0.09360263454777973   0.29121742621456825   0.10773753752104558
0.5196361990040789   0.6427332473608911   0.5120468644770008   0.926650655216808   0.23727357153143872   0.7771375013963113   0.7550527379344946   0.3585652175662597   0.3140041405903004   0.5129495451529847   0.6395827372055752   0.6300038525059257   0.7548864884890356   0.34694350825921244   0.5348396948547814   0.860772903052507   0.14752996317474332   0.7774683915425481   0.7673312010319121   0.4286570164803598   0.8251749166428032   0.6838657569947684   0.4761137748173438   0.3209194789593142   0.30553871763872426   0.041132509633877226   0.9640669103403431   0.39426882374250627   0.06826514610728551   0.2639950082375659   0.20901417240584846   0.0357036061762466   0.7542610055169852   0.7510454630845811   0.5694314352002733   0.40569975367032085   0.9993745170279495   0.40410195482536865   0.034591740345491874   0.5449268506178139   0.8518445538532062   0.6266335632828206   0.2672605393135798   0.11626983413745404   0.026669637210403094   0.9427678062880521   0.791146764496236   0.7953503551781398   0.7211309195716789   0.901635296654175   0.8270798541558929   0.4010815314356335   0.6528657734643933   0.637640288416609   0.6180656817500445   0.36537792525938695   0.8986047679474082   0.8865948253320279   0.0486342465497712   0.9596781715890661   0.8992302509194586   0.48249287050665934   0.014042506204279328   0.4147513209712522
0.04738569706625243   0.8558593072238387   0.7467819668906995   0.29848148683379816   0.02071605985584934   0.9130915009357866   0.9556352023944635   0.5031311316556584   0.2995851402841705   0.011456204281611652   0.12855534823857054   0.10204960022002482   0.6467193668197772   0.37381591586500257   0.5104896664885261   0.7366716749606379   0.748114598872369   0.4872210905329746   0.4618554199387549   0.7769935033715718   0.8488843479529102   0.00472822002631527   0.44781291373447557   0.36224218240031963   0.8014986508866578   0.1488689128024765   0.701030946843776   0.06376069556652145   0.7807825910308085   0.2357774118666899   0.7453957444493126   0.560629563910863   0.481197450746638   0.22432120758507826   0.6168403962107419   0.45857996369083825   0.8344780839268608   0.8505052917200757   0.1063507297222159   0.7219082887302004   0.08636348505449193   0.3632842011871011   0.644495309783461   0.9449147853586286   0.23747913710158167   0.3585559811607858   0.1966823960489855   0.5826726029583089   0.43598048621492386   0.2096870683583093   0.4956514492052095   0.5189119073917875   0.6551978951841154   0.9739096564916194   0.750255704755897   0.9582823434809244   0.1740004444374774   0.7495884489065412   0.13341530854515496   0.49970237979008614   0.3395223605106165   0.8990831571864655   0.02706457882293905   0.7777940910598857
0.2531588754561246   0.5357989559993644   0.382569269039478   0.8328793057012572   0.015679738354542935   0.17724297483857862   0.18588687299049253   0.2502067027429482   0.579699252139619   0.9675559064802693   0.690235423785283   0.7312947953511607   0.9245013569555037   0.9936462499886499   0.9399797190293862   0.7730124518702363   0.7505009125180263   0.24405780108210873   0.8065644104842312   0.2733100720801501   0.41097855200740974   0.34497464389564325   0.7794998316612921   0.4955159810202644   0.15781967655128515   0.8091756878962788   0.3969305626218141   0.6626366753190072   0.14213993819674223   0.6319327130577002   0.21104368963132158   0.412429972576059   0.5624406860571232   0.6643768065774309   0.5208082658460386   0.6811351772248982   0.6379393291016194   0.670730556588781   0.5808285468166524   0.908122725354662   0.8874384165835931   0.4266727555066723   0.7742641363324212   0.6348126532745119   0.4764598645761834   0.08169811161102902   0.9947643046711291   0.13929667225424747   0.31864018802489824   0.2725224237147502   0.5978337420493149   0.47665999693524025   0.17650024982815601   0.64058971065705   0.3867900524179934   0.06423002435918125   0.6140595637710329   0.9762129040796191   0.8659817865719549   0.383094847134283   0.9761202346694134   0.30548234749083814   0.2851532397553025   0.47497212177962095
0.08868181808582028   0.8788095919841659   0.5108891034228813   0.8401594685051091   0.6122219535096369   0.7971114803731368   0.5161247987517522   0.7008627962508617   0.29358176548473863   0.5245890566583866   0.9182910567024372   0.2242027993156214   0.11708151565658263   0.8839993460013367   0.5315010042844438   0.15997277495644013   0.5030219518855498   0.9077864419217175   0.6655192177124889   0.7768779278221571   0.5269017172161363   0.6023040944308794   0.38036597795718646   0.3019058060425362   0.43821989913031606   0.7234945024467135   0.8694768745343052   0.4617463375374271   0.8259979456206792   0.9263830220735767   0.35335207578255295   0.7608835412865654   0.5324161801359405   0.4017939654151901   0.4350610190801158   0.5366807419709441   0.4153346644793579   0.5177946194138534   0.9035600147956719   0.37670796701450393   0.9123127125938082   0.6100081774921359   0.23804079708318301   0.5998300391923468   0.3854109953776718   0.007704083061256495   0.8576748191259966   0.29792423314981054   0.9471910962473558   0.28420958061454293   0.9881979445916914   0.8361778956123834   0.12119315062667659   0.35782655854096623   0.6348458688091384   0.07529435432581798   0.5887769704907361   0.9560325931257762   0.19978484972902266   0.5386136123548739   0.17344230601137817   0.4382379737119227   0.2962248349333507   0.16190564534036997
0.26112959341757   0.8282297962197868   0.05818403785016767   0.5620756061480232   0.8757185980398982   0.8205257131585303   0.2005092187241711   0.2641513729982126   0.9285275017925424   0.5363161325439874   0.2123112741324797   0.4279734773858292   0.8073343511658658   0.17848957400302112   0.5774654053233412   0.3526791230600112   0.21855738067512978   0.222456980877245   0.3776805555943186   0.8140655107051373   0.04511507466375163   0.7842190071653223   0.0814557206609679   0.6521598653647673   0.7839854812461816   0.9559892109455356   0.023271682810800227   0.09008425921674414   0.9082668832062835   0.1354634977870053   0.8227624640866291   0.8259328862185314   0.979739381413741   0.599147365243018   0.6104511899541495   0.3979594088327023   0.17240503024787515   0.42065779123999686   0.032985784630808195   0.045280285772691116   0.9538476495727454   0.19820081036275186   0.6553052290364896   0.23121477506755383   0.9087325749089937   0.4139818031974295   0.5738495083755217   0.5790549097027865   0.12474709366281211   0.4579925922518939   0.5505778255647215   0.4889706504860424   0.21648021045652868   0.32252909446488864   0.7278153614780923   0.6630377642675108   0.2367408290427877   0.7233817292218706   0.11736417152394289   0.26507835543480857   0.06433579879491255   0.30272393798187375   0.08437838689313469   0.21979806966211743
0.1104881492221672   0.10452312761912191   0.42907315785664507   0.9885832945945636   0.20175557431317345   0.6905413244216924   0.8552236494811234   0.4095283848917771   0.07700848065036134   0.23254873216979843   0.30464582391640194   0.9205577344057347   0.8605282701938326   0.9100196377049098   0.5768304624383096   0.25751997013822386   0.623787441151045   0.18663790848303918   0.4594662909143667   0.9924416147034153   0.5594516423561324   0.8839139705011654   0.37508790402123204   0.772643545041298   0.4489634931339652   0.7793908428820435   0.9460147461645869   0.7840602504467343   0.24720791882079177   0.0888495184603511   0.09079109668346352   0.3745318655549572   0.1701994381704304   0.8563007862905527   0.7861452727670616   0.45397413114922247   0.30967116797659777   0.9462811485856428   0.209314810328752   0.19645416101099858   0.6858837268255528   0.7596432401026036   0.7498485194143852   0.20401254630758323   0.1264320844694204   0.8757292696014383   0.37476061539315325   0.4313690012662853   0.6774685913354552   0.0963384267193948   0.42874586922856633   0.647308750819551   0.43026067251466343   0.00748890825904369   0.3379547725451028   0.27277688526459376   0.260061234344233   0.15118812196849102   0.5518094997780412   0.8188027541153713   0.9503900663676352   0.20490697338284816   0.34249468944928924   0.6223485931043727
0.26450633954208247   0.44526373328024443   0.5926461700349039   0.4183360467967895   0.13807425507266208   0.5695344636788061   0.21788555464175072   0.9869670455305042   0.4606056637372069   0.47319603695941137   0.7891396854131844   0.3396582947109532   0.030344991222543475   0.4657071287003677   0.4511849128680816   0.06688140944635944   0.7702837568783104   0.31451900673187666   0.8993754130900404   0.2480786553309881   0.8198936905106752   0.10961203334902851   0.5568807236407511   0.6257300622266154   0.5553873509685927   0.6643483000687841   0.9642345536058472   0.20739401542982586   0.4173130958959307   0.09481383638997788   0.7463489989640965   0.22042696989932167   0.9567074321587238   0.6216177994305665   0.9572093135509121   0.8807686751883684   0.9263624409361803   0.15591067073019885   0.5060244006828305   0.813887265742009   0.15607868405786982   0.8413916639983222   0.6066489875927901   0.5658086104110209   0.3361849935471946   0.7317796306492936   0.04976826395203895   0.9400785481844055   0.7807976425786018   0.06743133058050964   0.08553371034619177   0.7326845327545797   0.3634845466826712   0.9726174941905318   0.3391847113820953   0.512257562855258   0.4067771145239475   0.35099969475996523   0.3819753978311832   0.6314888876668896   0.4804146735877672   0.19508902402976638   0.8759509971483528   0.8176016219248805
0.32433598952989734   0.3536973600314442   0.26930200955556266   0.25179301151385963   0.9881509959827027   0.6219177293821505   0.21953374560352373   0.3117144633294541   0.20735335340410083   0.5544863988016409   0.13400003525733195   0.5790299305748744   0.8438688067214296   0.5818689046111091   0.7948153238752367   0.06677236771961644   0.4370916921974821   0.23086920985114387   0.4128399260440534   0.4352834800527269   0.9566770186097149   0.0357801858213775   0.5368889288957006   0.6176818581278464   0.6323410290798176   0.6820828257899333   0.26758691934013795   0.36588884661398674   0.6441900330971149   0.060165096407782816   0.04805317373661425   0.054174383284532654   0.436836679693014   0.5056786976061419   0.9140531384792823   0.4751444527096582   0.5929678729715844   0.9238097929950329   0.11923781460404564   0.4083720849900418   0.15587618077410226   0.692940583143889   0.7063978885599922   0.9730886049373149   0.19919916216438735   0.6571603973225114   0.16950895966429158   0.35540674680946854   0.5668581330845698   0.9750775715325781   0.9019220403241536   0.9895179001954818   0.9226680999874549   0.9149124751247953   0.8538688665875394   0.9353435169109492   0.48583142029444093   0.40923377751865336   0.9398157281082571   0.4601990642012909   0.8928635473228566   0.4854239845236205   0.8205779135042114   0.051826979211249125
0.7369873665487543   0.7924834013797315   0.1141800249442192   0.07873837427393422   0.5377882043843669   0.1353230040572201   0.9446710652799276   0.7233316274644657   0.9709300712997971   0.16024543252464193   0.04274902495577401   0.7338137272689839   0.048261971312342236   0.24533295739984662   0.18888015836823466   0.7984702103580348   0.5624305510179013   0.8360991798811932   0.2490644302599776   0.33827114615674386   0.6695670036950447   0.3506751953575727   0.4284865167557662   0.28644416694549474   0.9325796371462904   0.5581917939778411   0.314306491811547   0.2077057926715605   0.3947914327619235   0.42286878992062105   0.3696354265316194   0.4843741652070948   0.4238613614621264   0.26262335739597914   0.32688640157584536   0.7505604379381109   0.37559939014978416   0.017290399996132525   0.1380062432076107   0.9520902275800761   0.8131688391318829   0.1811912201149393   0.8889418129476331   0.6138190814233323   0.14360183543683808   0.8305160247573666   0.4604552961918669   0.32737491447783756   0.2110221982905476   0.27232423077952544   0.1461488043803199   0.1196691218062771   0.8162307655286241   0.8494554408589043   0.7765133778487006   0.6352949565991823   0.3923694040664977   0.5868320834629253   0.4496269762728552   0.8847345186610714   0.016770013916713532   0.5695416834667927   0.31162073306524446   0.9326442910809952
0.2036011747848307   0.3883504633518534   0.4226789201176114   0.3188252096576629   0.059999339347992606   0.5578344385944868   0.9622236239257445   0.9914502951798253   0.848977141057445   0.2855102078149614   0.8160748195454245   0.8717811733735482   0.032746375528820953   0.43605476695605705   0.039561441696724   0.23648621677436596   0.6403769714623233   0.8492226834931318   0.5899344654238688   0.35175169811329454   0.6236069575456098   0.2796810000263391   0.27831373235862433   0.4191074070322993   0.42000578276077905   0.8913305366744857   0.855634812241013   0.10028219737463635   0.3600064434127864   0.33349609807999886   0.8934111883152686   0.108831902194811   0.5110293023553415   0.04798589026503746   0.07733636876984397   0.23705072882126274   0.4782829268265205   0.6119311233089805   0.03777492707311996   0.0005645120468967895   0.8379059553641972   0.7627084398158486   0.4478404616492511   0.6488128139336022   0.21429899781858747   0.4830274397895095   0.1695267292906268   0.22970540690130292   0.7942932150578084   0.5916969031150238   0.31389191704961383   0.12942320952666658   0.434286771645022   0.25820080503502496   0.42048072873434533   0.02059130733185558   0.9232574692896806   0.2102149147699875   0.3431443599645013   0.7835405785105929   0.44497454246316004   0.5982837914610071   0.3053694328913814   0.782976066463696
0.6070685870989628   0.8355753516451585   0.8575289712421302   0.1341632525300938   0.39276958928037536   0.35254791185564893   0.6880022419515035   0.9044578456287908   0.5984763742225669   0.7608510087406252   0.37411032490188967   0.7750346361021243   0.16418960257754495   0.5026502037056002   0.9536295961675443   0.7544433287702688   0.24093213328786442   0.2924352889356127   0.610485236203043   0.9709027502596759   0.7959575908247044   0.6941514974746057   0.3051158033116616   0.18792668379597985   0.18888900372574155   0.8585761458294472   0.44758683206953137   0.05376343126588602   0.7961194144453662   0.5060282339737983   0.7595845901180279   0.14930558563709515   0.19764304022279927   0.7451772252331731   0.38547426521613826   0.37427094953497086   0.03345343764525432   0.24252702152757294   0.4318446690485939   0.6198276207647021   0.7925213043573899   0.9500917325919602   0.8213594328455509   0.6489248705050262   0.9965637135326855   0.2559402351173546   0.5162436295338894   0.4609981867090464   0.8076747098069439   0.3973640892879074   0.06865679746435799   0.4072347554431604   0.011555295361577735   0.8913358553141091   0.3090722073463301   0.25792916980606523   0.8139122551387784   0.146158630080936   0.9235979421301919   0.8836582202710944   0.7804588174935242   0.9036316085533631   0.49175327308159794   0.26383059950639226
0.9879375131361342   0.9535398759614029   0.670393840236047   0.6149057290013661   0.9913737996034487   0.6975996408440482   0.15415021070215765   0.15390754229231965   0.1836990897965048   0.3002355515561409   0.08549341323779966   0.7466727868491593   0.17214379443492706   0.40889969624203176   0.7764212058914696   0.48874361704309405   0.3582315392961486   0.26274106616109577   0.8528232637612777   0.6050853967719997   0.5777727218026245   0.3591094576077327   0.3610699906796798   0.34125479726560737   0.5898352086664902   0.4055695816463299   0.6906761504436328   0.7263490682642413   0.5984614090630415   0.7079699408022816   0.5365259397414752   0.5724415259719217   0.41476231926653667   0.4077343892461407   0.45103252650367553   0.8257687391227624   0.24261852483160962   0.9988346930041089   0.674611320612206   0.33702512207966834   0.884386985535461   0.7360936268430132   0.8217880568509283   0.7319397253076687   0.30661426373283657   0.3769841692352804   0.46071806617124844   0.39068492804206134   0.7167790550663463   0.9714145875889505   0.7700419157276156   0.6643358597778201   0.11831764600330485   0.2634446467866689   0.23351597598614046   0.09189433380589834   0.7035553267367681   0.8557102575405282   0.782483449482465   0.26612559468313596   0.46093680190515857   0.8568755645364193   0.10787212887025897   0.9291004726034676
0.5765498163696976   0.12078193769340617   0.2860840720193307   0.19716074729579894   0.269935552636861   0.7437977684581257   0.8253660058480823   0.8064758192537376   0.5531564975705147   0.7723831808691752   0.05532409012046664   0.14213995947591762   0.4348388515672098   0.5089385340825063   0.8218081141343262   0.050245625670019264   0.7312835248304417   0.6532282765419781   0.039324664651861255   0.7841200309868833   0.27034672292528306   0.7963527120055589   0.9314525357816023   0.8550195583834157   0.6937969065555856   0.6755707743121527   0.6453684637622715   0.6578588110876168   0.42386135391872454   0.9317730058540269   0.8200024579141892   0.8513829918338791   0.8707048563482098   0.15938982498485166   0.7646783677937227   0.7092430323579615   0.435866004781   0.6504512909023453   0.9428702536593965   0.6589974066879423   0.7045824799505584   0.9972230143603672   0.9035455890075352   0.874877375701059   0.43423575702527534   0.2008703023548083   0.9720930532259329   0.019857817317643262   0.7404388504696898   0.5252995280426556   0.32672458946366134   0.3619990062300265   0.3165774965509653   0.5935265221886287   0.5067221315494721   0.5106160143961473   0.4458726402027554   0.434136697203777   0.7420437637557494   0.8013729820381859   0.010006635421755375   0.7836854063014317   0.799173510096353   0.14237557535024364
0.305424155471197   0.7864623919410645   0.8956279210888178   0.2674981996491847   0.8711883984459217   0.5855920895862562   0.9235348678628849   0.24764038233154143   0.13074954797623187   0.06029256154360066   0.5968102783992235   0.8856413761015149   0.8141720514252666   0.466766039354972   0.09008814684975147   0.3750253617053675   0.3682994112225112   0.032629342151195   0.34804438309400204   0.5736523796671816   0.3582927758007558   0.24894393584976332   0.548870872997649   0.431276804316938   0.05286862032955882   0.4624815439086988   0.6532429519088312   0.16377860466775332   0.18168022188363717   0.8768894543224426   0.7297080840459463   0.9161382223362119   0.05093067390740531   0.8165968927788418   0.13289780564672277   0.03049684623469698   0.23675862248213872   0.3498308534238699   0.0428096587969713   0.6554714845293295   0.8684592112596276   0.3172015112726749   0.6947652757029693   0.08181910486214786   0.5101664354588717   0.06825757542291157   0.14589440270532025   0.6505423005452099   0.45729781512931295   0.6057760315142128   0.49265145079648903   0.48676369587745655   0.27561759324567575   0.7288865771917703   0.7629433667505428   0.5706254735412447   0.22468691933827045   0.9122896844129283   0.6300455611038199   0.5401286273065476   0.9879282968561317   0.5624588309890585   0.5872359023068486   0.8846571427772182
0.11946908559650417   0.24525731971638362   0.8924706266038793   0.8028380379150704   0.6093026501376324   0.17699974429347204   0.7465762238985592   0.1522957373698605   0.15200483500831946   0.5712237127792592   0.2539247731020701   0.665532041492404   0.8763872417626437   0.842337135587489   0.49098140635152737   0.09490656795115929   0.6517003224243733   0.9300474511745607   0.8609358452477075   0.5547779406446116   0.6637720255682416   0.36758862018550215   0.2736999429408588   0.6701207978673934   0.5443029399717374   0.12233130046911851   0.3812293163369795   0.8672827599523231   0.9350002898341049   0.9453315561756465   0.6346530924384204   0.7149870225824626   0.7829954548257855   0.3741078433963872   0.38072831933635026   0.04945498109005861   0.9066082130631418   0.5317707078088982   0.8897469129848229   0.9545484131388993   0.2549078906387685   0.6017232566343376   0.028811067737115382   0.3997704724942877   0.591135865070527   0.23413463644883548   0.7551111247962565   0.7296496746268943   0.04683292509878964   0.11180333597971698   0.3738818084592771   0.8623669146745713   0.1118326352646847   0.16647177980407052   0.7392287160208567   0.14737989209210867   0.32883718043889926   0.7923639364076833   0.35850039668450645   0.09792491100205007   0.4222289673757575   0.2605932285987851   0.4687534836996836   0.14337649786315074
0.167321076736989   0.6588699719644474   0.4399424159625682   0.743606025368863   0.576185211666462   0.424735335515612   0.6848312911663117   0.013956350741968744   0.5293522865676724   0.312931999535895   0.3109494827070346   0.1515894360673975   0.4175196513029877   0.1464602197318245   0.5717207666861779   0.004209543975288827   0.08868247086408841   0.3540962833241412   0.21322037000167143   0.9062846329732388   0.6664535034883309   0.09350305472535614   0.7444668863019878   0.762908135110088   0.4991324267513419   0.4346330827609087   0.30452447033941954   0.019302109741224968   0.9229472150848799   0.009897747245296703   0.6196931791731078   0.0053457589992562254   0.3935949285172075   0.6969657477094017   0.30874369646607325   0.8537563229318588   0.9760752772142198   0.5505055279775772   0.7370229297798954   0.8495467789565699   0.8873928063501314   0.196409244653436   0.5238025597782239   0.9432621459833311   0.22093930286180052   0.10290618992807987   0.7793356734762361   0.18035401087324313   0.7218068761104586   0.6682731071671711   0.4748112031368166   0.16105190113201814   0.7988596610255787   0.6583753599218745   0.8551180239637087   0.15570614213276193   0.40526473250837125   0.9614096122124728   0.5463743274976355   0.3019498192009032   0.42918945529415137   0.41090408423489555   0.8093513977177401   0.4524030402443333
0.5417966489440199   0.21449483958145957   0.2855488379395162   0.5091408942610022   0.32085734608221944   0.1115886496533797   0.50621316446328   0.3287868833877591   0.5990504699717608   0.4433155424862085   0.03140196132646352   0.1677349822557409   0.800190808946182   0.7849401825643341   0.17628393736275483   0.012028840122978977   0.3949260764378108   0.8235305703518613   0.6299096098651193   0.7100790209220758   0.9657366211436594   0.4126264861169657   0.8205582121473793   0.25767598067774244   0.42393997219963947   0.1981316465355061   0.5350093742078631   0.7485350864167403   0.10308262611742008   0.0865429968821264   0.02879620974458305   0.4197482030289812   0.5040321561456593   0.6432274543959179   0.9973942484181195   0.2520132207732403   0.7038413471994772   0.8582872718315838   0.8211103110553647   0.23998438065026131   0.3089152707616664   0.03475670147972263   0.1912007011902453   0.5299053597281855   0.343178649618007   0.6221302153627569   0.37064248904286595   0.2722293790504431   0.9192386774183675   0.42399856882725084   0.8356331148350029   0.5236942926337028   0.8161560513009474   0.3374555719451245   0.8068369050904198   0.10394608960472164   0.3121238951552881   0.6942281175492065   0.8094426566723003   0.8519328688314813   0.6082825479558108   0.8359408457176227   0.9883323456169356   0.61194848818122
0.29936727719414447   0.8011841442379001   0.7971316444266903   0.08204312845303444   0.9561886275761374   0.17905392887514313   0.4264891553838243   0.8098137494025913   0.036949950157769994   0.7550553600478922   0.5908560405488215   0.2861194567688885   0.22079389885682257   0.41759978810276777   0.7840191354584016   0.18217336716416685   0.9086700037015345   0.7233716705535612   0.9745764787861014   0.33024049833268554   0.30038745574572356   0.8874308248359385   0.9862441331691658   0.7182920101514655   0.0010201785515791244   0.08624668059803839   0.1891124887424755   0.6362488816984311   0.04483155097544164   0.9071927517228953   0.7626233333586512   0.8264351322958398   0.00788160081767165   0.15213739167500304   0.1717672928098297   0.5403156755269513   0.7870877019608491   0.7345376035722353   0.38774815735142804   0.3581423083627844   0.8784176982593146   0.011165933018674072   0.41317167856532666   0.027901810030098874   0.578030242513591   0.1237351081827356   0.42692754539616085   0.30960979987863335   0.5770100639620119   0.03748842758469721   0.23781505665368535   0.6733609181802023   0.5321785129865703   0.13029567586180194   0.4751917232950342   0.8469257858843625   0.5242969121688986   0.978158284186799   0.3034244304852045   0.30661011035741126   0.7372092102080495   0.24362068061456366   0.9156762731337764   0.9484678019946269
0.8587915119487349   0.23245474759588958   0.5025045945684498   0.9205659919645279   0.2807612694351439   0.10871963941315398   0.07557704917228895   0.6109561920858946   0.703751205473132   0.07123121182845676   0.8377619925186036   0.9375952739056923   0.1715726924865618   0.9409355359666548   0.3625702692235694   0.09066948802132985   0.6472757803176632   0.962777251779856   0.059145838738364924   0.7840593776639186   0.9100665701096137   0.7191565711652923   0.14346956560458848   0.8355915756692918   0.05127505816087872   0.4867018235694027   0.6409649710361387   0.9150255837047637   0.7705137887257348   0.37798218415624874   0.5653879218638497   0.30406939161886914   0.06676258325260279   0.30675097232779197   0.7276259293452462   0.3664741177131768   0.895189890766041   0.36581543636113717   0.36505566012167673   0.27580462969184694   0.24791411044837783   0.4030381845812812   0.3059098213833118   0.49174525202792835   0.3378475403387642   0.683881613415989   0.1624402557787233   0.6561536763586366   0.28657248217788545   0.19717978984658624   0.5214752847425846   0.7411280926538728   0.5160586934521506   0.8191976056903375   0.956087362878735   0.4370587010350037   0.44929611019954785   0.5124466333625456   0.2284614335334888   0.07058458332182693   0.5541062194335069   0.1466311970014084   0.8634057734118121   0.79477995362998
0.30619210898512905   0.7435930124201272   0.5574959520285003   0.30303470160205165   0.9683445686463649   0.05971139900413821   0.395055696249777   0.6468810252434151   0.6817720864684794   0.862531609157552   0.8735804115071923   0.9057529325895423   0.16571339301632876   0.04333400346721446   0.9174930486284574   0.46869423155453854   0.7164172828167809   0.5308873701046689   0.6890316150949686   0.3981096482327116   0.16231106338327403   0.38425617310326055   0.8256258416831566   0.6033296946027316   0.856118954398145   0.6406631606831333   0.26812988965465623   0.3002949930006799   0.8877743857517801   0.5809517616789952   0.8730741934048792   0.6534139677572648   0.2060022992833007   0.7184201525214432   0.9994937818976869   0.7476610351677226   0.04028890626697194   0.6750861490542287   0.08200073326922949   0.2789668036131841   0.32387162345019105   0.14419877894955982   0.3929691181742609   0.8808571553804725   0.16156056006691702   0.7599426058462992   0.5673432764911044   0.2775274607777409   0.30544160566877204   0.11927944516316592   0.2992133868364481   0.977232467777061   0.4176672199169919   0.5383276834841707   0.42613919343156886   0.3238185000197961   0.21166492063369122   0.8199075309627276   0.42664541153388197   0.5761574648520735   0.1713760143667193   0.14482138190849883   0.34464467826465245   0.29719066123888943
0.8475043909165283   0.0006226029589389988   0.9516755600903916   0.41633350585841694   0.6859438308496112   0.2406799971126397   0.3843322835992872   0.1388060450806761   0.3805022251808392   0.12140055194947379   0.08511889676283911   0.16157357730361513   0.9628350052638472   0.583072868465303   0.6589797033312702   0.837755077283819   0.7511700846301561   0.7631653375025754   0.23233429179738826   0.2615976124317455   0.5797940702634368   0.6183439555940766   0.8876896135327358   0.964406951192856   0.7322896793469086   0.6177213526351376   0.9360140534423442   0.5480734453344391   0.046345848497297316   0.37704135552249796   0.551681769843057   0.409267400253763   0.6658436233164581   0.25564080357302416   0.4665628730802179   0.24769382295014788   0.7030086180526108   0.6725679351077212   0.8075831697489476   0.4099387456663289   0.9518385334224548   0.9094025976051456   0.5752488779515594   0.1483411332345834   0.372044463159018   0.291058642011069   0.6875592644188235   0.18393418204172737   0.6397547838121095   0.6733372893759314   0.7515452109764793   0.6358607367072883   0.5934089353148122   0.29629593385343345   0.19986344113342236   0.22659333645352528   0.927565311998354   0.0406551302804093   0.7333005680532044   0.9788995135033774   0.22455669394574318   0.3680871951726882   0.9257173983042568   0.5689607678370485
0.2727181605232884   0.45868459756754254   0.35046852035269743   0.4206196346024651   0.9006736973642704   0.1676259555564735   0.6629092559338738   0.23668545256073775   0.2609189135521609   0.4942886661805421   0.9113640449573945   0.6008247158534494   0.6675099782373488   0.19799273232710868   0.7115006038239721   0.3742313793999242   0.7399446662389947   0.15733760204669936   0.9782000357707676   0.3953318658965468   0.5153879722932515   0.7892504068740112   0.05248263746651084   0.8263710980594983   0.24266981176996313   0.33056580930646867   0.7020141171138135   0.40575146345703317   0.3419961144056928   0.16293985374999517   0.039104861179939575   0.16906601089629544   0.08107720085353184   0.6686511875694531   0.1277408162225451   0.5682412950428459   0.41356722261618306   0.4706584552423444   0.41624021239857295   0.1940099156429218   0.6736225563771884   0.313320853195645   0.4380401766278053   0.798678049746375   0.15823458408393684   0.5240704463216338   0.3855575391612945   0.9723069516868768   0.9155647723139737   0.19350463701516518   0.6835434220474811   0.5665554882298436   0.5735686579082809   0.03056478326517   0.6444385608675415   0.3974894773335481   0.49249145705474906   0.36191359569571696   0.5166977446449964   0.8292481822907022   0.078924234438566   0.8912551404533725   0.10045753224642343   0.6352382666477804
0.4053016780613776   0.5779342872577276   0.6624173556186181   0.8365602169014054   0.2470670939774408   0.05386384093609365   0.2768598164573236   0.8642532652145286   0.3315023216634671   0.8603592039209285   0.5933163944098425   0.2976977769846851   0.7579336637551862   0.8297944206557585   0.948877833542301   0.9002082996511369   0.2654422067004371   0.4678808249600415   0.4321800888973047   0.07096011736043482   0.1865179722618711   0.576625684506669   0.33172255665088124   0.43572185071265446   0.7812162942004934   0.9986913972489415   0.6693052010322631   0.5991616338112491   0.5341492002230527   0.9448275563128479   0.39244538457493955   0.7349083685967205   0.20264687855958555   0.08446835239191938   0.799128990165097   0.43721059161203546   0.44471321480439935   0.25467393173616093   0.8502511566227959   0.5370022919608984   0.17927100810396226   0.7867931067761194   0.41807106772549124   0.46604217460046365   0.9927530358420912   0.21016742226945037   0.08634851107460996   0.03032032388780918   0.2115367416415977   0.21147602502050886   0.4170433100423468   0.43115869007656005   0.6773875414185451   0.266648468707661   0.024597925467407283   0.6962503214798396   0.47474066285895944   0.18218011631574163   0.22546893530231032   0.2590397298678041   0.0300274480545601   0.9275061845795807   0.37521777867951445   0.7220374379069057
0.8507564399505978   0.14071307780346134   0.9571467109540231   0.25599526330644196   0.8580034041085067   0.930545655534011   0.8707981998794132   0.2256749394186328   0.646466662466909   0.7190696305135021   0.4537548898370664   0.7945162493420728   0.969079121048364   0.45242116180584113   0.42915696436965917   0.0982659278622332   0.49433845818940453   0.27024104549009953   0.2036880290673488   0.8392261979944291   0.4643110101348444   0.3427348609105188   0.8284702503878344   0.11718876008752345   0.6135545701842465   0.20202178310705746   0.8713235394338112   0.8611934967810815   0.7555511660757399   0.27147612757304646   0.000525339554397968   0.6355185573624487   0.1090845036088309   0.5524064970595444   0.5467704497173316   0.8410023080203759   0.14000538256046693   0.09998533525370322   0.1176134853476724   0.7427363801581427   0.6456669243710624   0.8297442897636037   0.9139254562803236   0.9035101821637136   0.18135591423621802   0.4870094288530849   0.08545520589248917   0.7863214220761902   0.5678013440519715   0.2849876457460275   0.21413166645867796   0.9251279252951087   0.8122501779762316   0.013511518172980982   0.21360632690428   0.28960936793266   0.7031656743674006   0.46110502111343665   0.6668358771869485   0.4486070599122841   0.5631602918069337   0.3611196858597334   0.549222391839276   0.7058706797541414
0.9174933674358713   0.5313753960961297   0.6352969355589525   0.8023604975904277   0.7361374531996533   0.04436596724304482   0.5498417296664633   0.01603907551423756   0.16833610914768188   0.7593783214970173   0.33571006320778535   0.09091115021912885   0.3560859311714503   0.7458668033240364   0.12210373630350536   0.8013017822864689   0.6529202568040496   0.2847617822105997   0.4552678591165569   0.3526947223741847   0.0897599649971159   0.9236420963508664   0.9060454672772809   0.6468240426200433   0.17226659756124457   0.3922667002547366   0.27074853171832836   0.8444635450296156   0.4361291443615913   0.3479007330116918   0.7209068020518651   0.8284244695153781   0.2677930352139094   0.5885224115146744   0.38519673884407973   0.7375133192962492   0.9117071040424591   0.842655608190638   0.2630930025405744   0.9362115370097803   0.25878684723840945   0.5578938259800382   0.8078251434240175   0.5835168146355957   0.16902688224129353   0.634251729629172   0.9017796761467366   0.9366927720155523   0.996760284680049   0.24198502937443536   0.6310311444284082   0.0922292269859367   0.5606311403184577   0.8940842963627436   0.9101243423765432   0.26380475747055865   0.2928381051045483   0.3055618848480692   0.5249276035324634   0.5262914381743095   0.3811310010620892   0.46290627665743117   0.26183460099188904   0.5900799011645291
0.12234415382367975   0.9050124506773929   0.4540094575678716   0.006563086528933444   0.9533172715823862   0.27076072104822096   0.552229781421135   0.06987031451338113   0.9565569869023373   0.028775691673785565   0.9211986369927267   0.9776410875274444   0.3959258465838796   0.13469139531104196   0.011074294616183653   0.7138363300568857   0.10308774147933127   0.8291295104629728   0.4861466910837202   0.1875448918825763   0.7219567404172421   0.36622323380554156   0.22431209009183117   0.5974649907180472   0.5996125865935623   0.46121078312814867   0.7703026325239596   0.5909019041891137   0.6462953150111761   0.19045006207992773   0.21807285110282457   0.5210315896757326   0.6897383281088388   0.16167437040614216   0.2968742141100978   0.5433905021482882   0.2938124815249593   0.026982975095100212   0.2857999194939141   0.8295541720914025   0.19072474004562803   0.19785346463212744   0.7996532284101939   0.6420092802088261   0.46876799962838595   0.8316302308265858   0.5753411383183628   0.044544289490778925   0.8691554130348237   0.3704194476984372   0.8050385057944032   0.4536423853016652   0.22286009802364756   0.17996938561850948   0.5869656546915786   0.9326107956259325   0.5331217699148088   0.018295015212367288   0.2900914405814808   0.38922029347764436   0.2393092883898494   0.991312040117267   0.004291521087566696   0.5596661213862419
0.04858454834422139   0.7934585754851396   0.20463829267737282   0.9176568411774157   0.5798165487158354   0.9618283446585537   0.6292971543590101   0.8731125516866368   0.7106611356810117   0.5914088969601166   0.824258648564607   0.4194701663849717   0.4878010376573642   0.4114395113416071   0.2372929938730284   0.4868593707590391   0.9546792677425555   0.3931444961292398   0.9472015532915475   0.0976390772813948   0.7153699793527061   0.4018324560119727   0.9429100322039808   0.5379729558951529   0.6667854310084848   0.608373880526833   0.7382717395266081   0.6203161147177371   0.08696888229264928   0.6465455358682793   0.10897458516759796   0.7472035630311002   0.3763077466116375   0.055136638908162804   0.284715936602991   0.3277333966461285   0.8885067089542733   0.6436971275665557   0.0474229427299626   0.8408740258870894   0.9338274412117178   0.25055263143731593   0.10022138943841502   0.7432349486056946   0.2184574618590117   0.8487201754253432   0.15731135723443412   0.2052619927105417   0.551672030850527   0.24034629489851012   0.41903961770782605   0.5849458779928046   0.4647031485578777   0.5938007590302308   0.3100650325402281   0.8377423149617044   0.08839540194624022   0.538664120122068   0.025349095937237085   0.5100089183155759   0.19988869299196693   0.8949669925555123   0.9779261532072745   0.6691348924284866
0.26606125178024914   0.6444143611181963   0.8777047637688594   0.925899943822792   0.04760378992123747   0.7956941856928531   0.7203934065344253   0.7206379511122503   0.49593175907071047   0.555347890794343   0.3013537888265993   0.13569207311944562   0.031228610512832752   0.9615471317641122   0.9912887562863713   0.2979497581577412   0.9428332085665926   0.4228830116420443   0.9659396603491341   0.7879408398421653   0.7429445155746256   0.5279160190865321   0.9880135071418596   0.1188059474136788   0.47688326379437646   0.8835016579683358   0.11030874337300017   0.19290600359088686   0.429279473873139   0.08780747227548268   0.3899153368385748   0.4722680524786366   0.9333477148024285   0.5324595814811397   0.08856154801197554   0.336575979359191   0.9021191042895957   0.5709124497170275   0.09727279172560432   0.03862622120144978   0.9592858957230032   0.14802943807498317   0.1313331313764702   0.2506853813592845   0.21634138014837762   0.6201134189884511   0.14331962423461056   0.13187943394560567   0.7394581163540012   0.7366117610201154   0.033010880861610394   0.9389734303547188   0.3101786424808622   0.6488042887446327   0.6430955440230356   0.46670537787608224   0.3768309276784337   0.11634470726349298   0.55453399601106   0.13012939851689123   0.47471182338883794   0.5454322575464655   0.4572612042854557   0.09150317731544146
0.5154259276658347   0.39740281947148237   0.3259280729089855   0.840817795956157   0.2990845475174571   0.7772894004830313   0.18260844867437492   0.7089383620105513   0.559626431163456   0.040677639462915936   0.14959756781276454   0.7699649316558325   0.24944778868259376   0.3918733507182833   0.506502023789729   0.3032595537797503   0.87261686100416   0.2755286434547903   0.951968027778669   0.17313015526285902   0.3979050376153221   0.7300963859083247   0.49470682349321327   0.08162697794741756   0.8824791099494873   0.3326935664368424   0.16877875058422775   0.24080918199126058   0.5833945624320303   0.5554041659538111   0.9861703019098528   0.5318708199807093   0.02376813126857425   0.5147265264908951   0.8365727340970883   0.7619058883248768   0.7743203425859805   0.1228531757726119   0.3300707103073593   0.45864633454512654   0.9017034815818205   0.8473245323178216   0.3781026825286904   0.2855161792822675   0.5037984439664983   0.11722814640949686   0.8833958590354771   0.20388920133484995   0.621319334017011   0.7845345799726545   0.7146171084512494   0.9630800193435893   0.03792477158498082   0.22913041401884335   0.7284468065413965   0.4312091993628801   0.014156640316406567   0.7144038875279481   0.8918740724443083   0.6693033110380033   0.23983629773042608   0.5915507117553362   0.5618033621369489   0.2106569764928768
0.33813281614860563   0.7442261794375147   0.18370067960825856   0.9251407972106093   0.8343343721821073   0.6269980330280178   0.3003048205727814   0.7212515958757594   0.21301503816509623   0.8424634530553633   0.585687712121532   0.7581715765321699   0.17509026658011542   0.61333303903652   0.8572409055801355   0.3269623771692899   0.16093362626370886   0.8989291515085718   0.9653668331358273   0.6576590661312866   0.9210973285332827   0.30737843975323553   0.40356347099887835   0.44700208963840976   0.5829645123846772   0.5631522603157209   0.2198627913906198   0.5218612924278004   0.7486301402025699   0.936154227287703   0.9195579708178384   0.8006096965520411   0.5356151020374736   0.09369077423233968   0.3338702586963063   0.042438120019871135   0.36052483545735825   0.4803577351958197   0.4766293531161708   0.7154757428505812   0.1995912091936494   0.5814285836872479   0.5112625199803436   0.05781667671929472   0.2784938806603666   0.2740501439340124   0.10769904898146516   0.610814587080885   0.6955293682756895   0.7108978836182915   0.8878362575908454   0.08895329465308452   0.9468992280731195   0.7747436563305885   0.968278286773007   0.28834359810104343   0.4112841260356459   0.6810528820982489   0.6344080280767007   0.24590547808117227   0.05075929057828765   0.20069514690242915   0.15777867496052994   0.530429735230591
0.8511680813846383   0.6192665632151813   0.6465161549801864   0.47261305851129626   0.5726742007242717   0.34521641928116886   0.5388171059987212   0.8617984714304113   0.8771448324485822   0.6343185356628773   0.650980848407876   0.7728451767773268   0.9302456043754627   0.8595748793322888   0.6827025616348689   0.4845015786762834   0.5189614783398168   0.17852199723403997   0.04829453355816817   0.23859610059511113   0.4682021877615291   0.9778268503316109   0.8905158585976383   0.7081663653645202   0.6170341063768908   0.3585602871164296   0.2439997036174518   0.23555330685322384   0.044359905652619186   0.01334386783526074   0.7051825976187305   0.3737548354228125   0.16721507320403697   0.37902533217238343   0.054201749210854626   0.6009096586454857   0.23696946882857434   0.5194504528400946   0.3714991875759857   0.11640807996920234   0.7180079904887575   0.3409284556060546   0.32320465401781756   0.8778119793740912   0.24980580272722847   0.3631016052744438   0.43268879542017935   0.1696456140095711   0.6327716963503376   0.004541318158014188   0.18868909180272753   0.9340923071563473   0.5884117906977184   0.9911974503227534   0.483506494183997   0.5603374717335348   0.4211967174936814   0.61217211815037   0.42930474497314236   0.959427813088049   0.18422724866510712   0.09272166531027543   0.05780555739715663   0.8430197331188466
0.46621925817634957   0.7517932097042208   0.734600903379339   0.9652077537447554   0.21641345544912108   0.388691604429777   0.30191210795915974   0.7955621397351843   0.5836417590987835   0.38415028627176284   0.11322301615643222   0.8614698325788371   0.995229968401065   0.39295283594900937   0.6297165219724352   0.30113236084530237   0.5740332509073837   0.7807807177986393   0.20041177699929286   0.3417045477572534   0.3898060022422765   0.688059052488364   0.14260621960213624   0.49868481463840675   0.9235867440659269   0.9362658427841432   0.4080053162227972   0.5334770608936513   0.7071732886168058   0.5475742383543661   0.10609320826363743   0.737914921158467   0.12353152951802238   0.1634239520826033   0.9928701921072052   0.8764450885796299   0.1283015611169573   0.770471116133594   0.36315367013476996   0.5753127277343275   0.5542683102095737   0.9896903983349546   0.16274189313547713   0.23360817997707412   0.16446230796729722   0.3016313458465907   0.02013567353334089   0.7349233653386674   0.24087556390137027   0.3653655030624476   0.6121303573105438   0.20144630444501607   0.5337022752845644   0.8177912647080814   0.5060371490469063   0.46353138328654914   0.41017074576654206   0.6543673126254781   0.513166956939701   0.5870862947069192   0.2818691846495847   0.8838961964918842   0.15001328680493112   0.011773566972591723
0.727600874440011   0.8942057981569296   0.987271393669454   0.7781653869955176   0.5631385664727138   0.5925744523103389   0.9671357201361132   0.04324202165685021   0.32226300257134355   0.22720894924789134   0.3550053628255694   0.8417957172118341   0.7885607272867791   0.4094176845398099   0.848968213778663   0.378264333925285   0.37838998152023706   0.7550503719143318   0.335801256838962   0.7911780392183658   0.09652079687065232   0.8711541754224476   0.18578797003403086   0.779404472245774   0.3689199224306413   0.976948377265518   0.19851657636457687   0.0012390852502564692   0.8057813559579274   0.3843739249551791   0.23138085622846377   0.9579970635934063   0.48351835338658394   0.15716497570728777   0.8763754934028944   0.11620134638157212   0.6949576260998048   0.7477472911674778   0.02740727962423132   0.7379370124562871   0.3165676445795678   0.9926969192531461   0.6916060227852693   0.9467589732379214   0.2200468477089155   0.12154274383069846   0.5058180527512385   0.16735450099214724   0.8511269252782742   0.14459436656518046   0.3073014763866616   0.16611541574189076   0.04534556932034672   0.7602204416100014   0.07592062015819781   0.2081183521484845   0.5618272159337627   0.6030554659027136   0.19954512675530342   0.09191700576691239   0.8668695898339579   0.8553081747352358   0.1721378471310721   0.3539799933106253
0.5503019452543901   0.8626112554820897   0.48053182434580277   0.407221020072704   0.3302550975454746   0.7410685116513912   0.9747137715945643   0.23986651908055676   0.4791281722672004   0.5964741450862108   0.6674122952079027   0.07375110333866598   0.43378260294685367   0.8362537034762094   0.5914916750497049   0.8656327511901815   0.8719553870130909   0.2331982375734958   0.39194654829440145   0.773715745423269   0.0050857971791330205   0.37789006283826004   0.21980870116332937   0.4197357521126438   0.4547838519247429   0.5152788073561704   0.7392768768175266   0.012514732039939799   0.1245287543792683   0.7742102957047792   0.7645631052229623   0.772648212959383   0.6454005821120679   0.1777361506185684   0.0971508100150596   0.698897109620717   0.21161797916521422   0.341482447142359   0.5056591349653548   0.8332643584305356   0.3396625921521233   0.1082842095688632   0.11371258667095323   0.05954861300726652   0.33457679497299025   0.7303941467306031   0.8939038855076239   0.6398128608946227   0.8797929430482473   0.21511533937443278   0.15462700869009727   0.627298128854683   0.755264188668979   0.4409050436696536   0.39006390346713493   0.8546499158952999   0.10986360655691113   0.2631688930510852   0.2929130934520754   0.15575280627458282   0.8982456273916969   0.9216864459087263   0.7872539584867206   0.32248844784404723
0.5585830352395736   0.8134022363398631   0.6735413718157675   0.2629398348367807   0.2240062402665834   0.0830080896092599   0.7796374863081436   0.623126973942158   0.34421329721833605   0.8678927502348271   0.6250104776180463   0.995828845087475   0.588949108549357   0.4269877065651735   0.23494657415091133   0.14117892919217515   0.4790855019924459   0.16381881351408828   0.942033480698836   0.9854261229175924   0.5808398746007489   0.24213236760536203   0.15477952221211533   0.6629376750735451   0.0222568393611753   0.428730131265499   0.4812381503963479   0.39999784023676443   0.798250599094592   0.3457220416562391   0.7016006640882043   0.7768708662946064   0.4540373018762559   0.477829291421412   0.07659018647015803   0.7810420212071314   0.8650881933268989   0.05084158485623849   0.8416436123192467   0.6398630920149563   0.38600269133445303   0.8870227713421502   0.8996101316204107   0.6544369690973639   0.805162816733704   0.6448904037367882   0.7448306094082954   0.9914992940238189   0.7829059773725288   0.2161602724712892   0.2635924590119475   0.5915014537870544   0.9846553782779368   0.8704382308150501   0.5619917949237432   0.814630587492448   0.530618076401681   0.3926089393936381   0.48540160845358515   0.03358856628531658   0.6655298830747821   0.3417673545373996   0.6437579961343385   0.3937254742703603
0.2795271917403291   0.4547445831952494   0.7441478645139278   0.7392885051729963   0.474364375006625   0.8098541794584612   0.9993172551056323   0.7477892111491774   0.6914583976340962   0.593693906987172   0.7357247960936848   0.15628775736212294   0.7068030193561594   0.7232556761721219   0.17373300116994164   0.3416571698696749   0.1761849429544784   0.33064673677848383   0.6883313927163565   0.30806860358435834   0.5106550598796963   0.9888793822410842   0.04457339658201805   0.9143431293139981   0.23112786813936723   0.5341347990458348   0.3004255320680903   0.17505462414100176   0.7567634931327423   0.7242806195873737   0.301108276962458   0.42726541299182436   0.06530509549864599   0.13058671260020163   0.5653834808687732   0.2709776556297014   0.35850207614248664   0.4073310364280797   0.39165047969883154   0.9293204857600265   0.18231713318800824   0.0766842996495959   0.703319086982475   0.6212518821756681   0.671662073308312   0.08780491740851169   0.6587456904004569   0.7069087528616701   0.4405342051689447   0.5536701183626769   0.35832015833236663   0.5318541287206683   0.6837707120362025   0.8293894987753032   0.05721188136990866   0.10458871572884394   0.6184656165375565   0.6988027861751016   0.4918284005011355   0.8336110600991425   0.25996354039506986   0.29147174974702184   0.10017792080230398   0.9042905743391161
0.07764640720706163   0.21478745009742595   0.39685883381982895   0.28303869216344796   0.4059843338987497   0.12698253268891427   0.738113143419372   0.5761299393017779   0.965450128729805   0.5733124143262374   0.3797929850870053   0.044275810581109604   0.2816794166936025   0.7439229155509341   0.3225811037170967   0.9396870948522656   0.663213800156046   0.0451201293758326   0.8307527032159612   0.10607603475312312   0.4032502597609761   0.7536483796288107   0.7305747824136573   0.20178546041400705   0.3256038525539145   0.5388609295313848   0.33371594859382825   0.9187467682505591   0.9196195186551648   0.4118783968424705   0.5956028051744563   0.3426168289487812   0.9541693899253598   0.8385659825162332   0.21580982008745092   0.29834101836767163   0.6724899732317573   0.09464306696529894   0.8932287163703543   0.3586539235154059   0.009276173075711288   0.04952293758946634   0.06247601315439307   0.2525778887622828   0.6060259133147352   0.2958745579606556   0.33190123074073585   0.050792428348275756   0.28042206076082066   0.7570136284292708   0.9981852821469076   0.13204566009771665   0.3608025421056559   0.34513523158680026   0.40258247697245136   0.7894288311489355   0.4066331521802961   0.5065692490705672   0.18677265688500044   0.49108781278126384   0.7341431789485388   0.4119261821052682   0.29354394051464616   0.1324338892658579
0.7248670058728275   0.3624032445158019   0.2310679273602531   0.879856000503575   0.11884109255809235   0.0665286865551463   0.8991666966195172   0.8290635721552994   0.8384190317972717   0.3095150581258755   0.9009814144726096   0.6970179120575827   0.4776164896916158   0.9643798265390752   0.49839893750015823   0.9075890809086472   0.07098333751131972   0.45781057746850806   0.31162628061515785   0.4165012681273834   0.33684015856278093   0.04588439536323981   0.018082340100511653   0.2840673788615255   0.6119731526899534   0.6834811508474379   0.7870144127402585   0.4042113783579504   0.49313206013186106   0.6169524642922917   0.8878477161207413   0.575147806202651   0.6547130283345894   0.3074374061664161   0.9868663016481317   0.8781298941450685   0.1770965386429736   0.34305757962734096   0.4884673641479734   0.9705408132364212   0.10611320113165387   0.8852470021588329   0.1768410835328156   0.5540395451090379   0.769273042568873   0.839362606795593   0.15875874343230395   0.2699721662475123   0.15729988987891952   0.15588145594815517   0.3717443306920454   0.8657607878895619   0.6641678297470585   0.5389289916558635   0.4838966145713041   0.2906129816869108   0.009454801412469039   0.2314915854894474   0.4970303129231724   0.4124830875418424   0.8323582627694954   0.8884340058621064   0.008562948775198974   0.44194227430542116
0.7262450616378415   0.003187003703273566   0.8317218652423833   0.8879027291963834   0.9569720190689687   0.16382439690768047   0.6729631218100794   0.617930562948871   0.7996721291900492   0.007942940959525309   0.301218791118034   0.7521697750593092   0.13550429944299067   0.46901394930366175   0.8173221765467299   0.46155679337239836   0.12604949803052165   0.23752236381421435   0.32029186362355755   0.049073705830556015   0.2936912352610262   0.3490883579521079   0.3117289148483586   0.6071314315251348   0.5674461736231846   0.34590135424883434   0.4800070496059752   0.7192287023287515   0.6104741545542159   0.18207695734115384   0.8070439277958957   0.10129813937988041   0.8108020253641669   0.17413401638162854   0.5058251366778618   0.34912836432057126   0.6752977259211762   0.7051200670779668   0.6885029601311318   0.8875715709481728   0.5492482278906545   0.46759770326375244   0.3682110965075742   0.8384978651176168   0.2555569926296284   0.11850934531164452   0.05648218165921567   0.231366433592482   0.6881108190064438   0.7726079910628102   0.5764751320532405   0.5121377312637305   0.07763666445222776   0.5905310337216564   0.7694312042573447   0.4108395918838501   0.2668346390880609   0.4163970173400278   0.263606067579483   0.06171122756327887   0.5915369131668847   0.7112769502620611   0.5751031074483512   0.17413965661510603
0.042288685276230135   0.2436792469983086   0.206892010940777   0.3356417914974892   0.7867316926466018   0.1251699016866641   0.15040982928156132   0.10427535790500718   0.09862087364015802   0.3525619106238539   0.5739346972283208   0.5921376266412767   0.020984209187930262   0.7620308769021975   0.8045034929709761   0.18129803475742656   0.7541495700998694   0.34563385956216974   0.5408974253914931   0.11958680719414767   0.16261265693298468   0.6343569093001087   0.9657943179431419   0.9454471505790417   0.12032397165675456   0.3906776623018001   0.7589023070023649   0.6098053590815525   0.33359227901015276   0.26550776061513603   0.6084924777208036   0.5055300011765453   0.23497140536999475   0.9129458499912821   0.03455778049248274   0.9133923745352687   0.2139871961820645   0.1509149730890846   0.2300542875215066   0.7320943397778421   0.45983762608219514   0.8052811135269149   0.6891568621300135   0.6125075325836944   0.2972249691492104   0.17092420422680613   0.7233625441868716   0.6670603820046528   0.17690099749245589   0.780246541925006   0.9644602371845067   0.057255022923100266   0.8433087184823032   0.5147387813098699   0.3559677594637032   0.5517250217465549   0.6083373131123083   0.6017929313185878   0.3214099789712204   0.6383326472112864   0.39435011693024385   0.45087795822950316   0.09135569144971381   0.9062383074334442
0.9345124908480487   0.6455968447025883   0.4021988293197003   0.2937307748497498   0.6372875216988383   0.47467264047578217   0.6788362851328287   0.6266703928450971   0.4603865242063824   0.6944260985507762   0.7143760479483219   0.5694153699219968   0.6170778057240793   0.17968731724090622   0.35840828848461875   0.017690348175441826   0.008740492611770949   0.5778943859223185   0.03699830951339832   0.3793577009641555   0.6143903756815271   0.12701642769281524   0.9456426180636845   0.4731193935307113   0.6798778848334784   0.4814195829902269   0.5434437887439842   0.17938861868096148   0.04259036313464013   0.006746942514444737   0.8646075036111556   0.5527182258358644   0.5822038389282578   0.31232084396366855   0.15023145566283366   0.9833028559138677   0.9651260332041784   0.13263352672276232   0.7918231671782149   0.9656125077384258   0.9563855405924075   0.5547391408004438   0.7548248576648166   0.5862548067742703   0.3419951649108804   0.42772271310762866   0.8091822396011321   0.11313541324355902   0.662117280077402   0.9463031301174017   0.26573845085714787   0.9337467945625976   0.6195269169427619   0.939556187602957   0.4011309472459923   0.38102856872673313   0.037323078014504116   0.6272353436392885   0.2508994915831586   0.39772571281286545   0.07219704481032566   0.4946018169165261   0.4590763244049437   0.4321132050744397
0.11581150421791814   0.9398626761160822   0.7042514667401272   0.8458583983001694   0.7738163393070377   0.5121399630084535   0.8950692271389951   0.7327229850566104   0.11169905922963573   0.5658368328910519   0.6293307762818472   0.7989761904940128   0.4921721422868739   0.6262806452880949   0.22819982903585492   0.4179476217672797   0.45484906427236976   0.9990453016488064   0.9773003374526963   0.02022190895441421   0.3826520194620441   0.5044434847322804   0.5182240130477526   0.5881087038799746   0.266840515244126   0.5645808086161982   0.8139725463076255   0.7422503055798052   0.49302417593708825   0.0524408456077446   0.9189033191686304   0.009527320523194863   0.3813251167074525   0.48660401271669274   0.2895725428867832   0.21055113002918208   0.8891529744205786   0.8603233674285978   0.061372713850928254   0.7926035082619024   0.4343039101482089   0.8612780657797914   0.08407237639823194   0.7723815993074882   0.051651890686164784   0.3568345810475109   0.5658483633504794   0.18427289542751363   0.7848113754420388   0.7922537724313128   0.7518758170428539   0.4420225898477084   0.2917871995049506   0.7398129268235681   0.8329724978742234   0.43249526932451354   0.9104620827974981   0.25320891410687546   0.5433999549874403   0.2219441392953315   0.021309108376919413   0.39288554667827763   0.4820272411365121   0.4293406310334291
0.5870051982287106   0.5316074808984863   0.3979548647382801   0.656959031725941   0.5353533075425457   0.17477289985097538   0.8321065013878007   0.4726861362984273   0.7505419321005069   0.3825191274196626   0.08023068434494687   0.0306635464507189   0.4587547325955564   0.6427062005960944   0.2472581864707234   0.5981682771262053   0.5482926497980583   0.389497286489219   0.7038582314832831   0.37622413783087383   0.5269835414211389   0.9966117398109414   0.22183099034677103   0.9468835067974447   0.9399783431924283   0.46500425891245506   0.8238761256084909   0.2899244750715038   0.4046250356498826   0.2902313590614797   0.9917696242206901   0.8172383387730765   0.6540831035493757   0.907712231641817   0.9115389398757433   0.7865747923223576   0.19532837095381936   0.2650060310457226   0.6642807534050199   0.18840651519615223   0.647035721155761   0.8755087445565036   0.9604225219217368   0.8121823773652784   0.12005217973462215   0.8788970047455622   0.7385915315749658   0.8652988705678336   0.18007383654219378   0.4138927458331072   0.9147154059664748   0.5753743954963298   0.7754488008923112   0.12366138677162751   0.9229457817457847   0.7581360567232533   0.12136569734293544   0.21594915512981042   0.011406841870041444   0.9715612644008957   0.9260373263891161   0.9509431240840878   0.3471260884650216   0.7831547492047436
0.27900160523335504   0.07543437952758417   0.38670356654328475   0.9709723718394652   0.1589494254987329   0.1965373747820219   0.6481120349683189   0.1056735012716315   0.9788755889565391   0.7826446289489147   0.7333966290018441   0.5302991057753017   0.20342678806422798   0.6589832421772872   0.8104508472560593   0.7721630490520482   0.08206109072129253   0.44303408704747677   0.7990440053860179   0.8006017846511525   0.15602376433217643   0.492090962963389   0.45191791692099637   0.01744703544640895   0.8770221590988214   0.4166565834358048   0.06521435037771162   0.0464746636069438   0.7180727336000885   0.2201192086537829   0.4171023154093927   0.9408011623353123   0.7391971446435494   0.4374745797048682   0.6837056864075486   0.41050205656001065   0.5357703565793214   0.778491337527581   0.8732548391514893   0.6383390075079624   0.45370926585802884   0.3354572504801042   0.07421083376547134   0.8377372228568098   0.2976855015258524   0.8433662875167152   0.622292916844475   0.8202901874104009   0.420663342427031   0.4267097040809104   0.5570785664667633   0.7738155238034571   0.7025906088269426   0.20659049542712749   0.1399762510573707   0.8330143614681448   0.9633934641833932   0.7691159157222593   0.4562705646498221   0.4225123049081342   0.4276231076040718   0.9906245781946783   0.5830157254983328   0.7841732974001718
0.973913841746043   0.6551673277145741   0.5088048917328615   0.946436074543362   0.6762283402201906   0.8118010401978589   0.8865119748883865   0.12614588713296102   0.25556499779315955   0.3850913361169485   0.32943340842162316   0.3523303633295039   0.552974388966217   0.178500840689821   0.18945715736425248   0.5193160018613591   0.5895809247828239   0.4093849249675617   0.7331865927144304   0.0968036969532249   0.161957817178752   0.4187603467728834   0.15017086721609757   0.3126303995530531   0.188043975432709   0.7635930190583092   0.641365975483236   0.3661943250096911   0.5118156352125185   0.9517919788604504   0.7548540005948495   0.2400484378767301   0.2562506374193589   0.5667006427435018   0.42542059217322636   0.8877180745472262   0.7032762484531419   0.3881998020536809   0.2359634348089739   0.36840207268586717   0.11369532367031808   0.9788148770861191   0.5027768420945435   0.2715983757326423   0.9517375064915661   0.5600545303132358   0.3526059748784459   0.9589679761795892   0.7636935310588571   0.7964615112549265   0.7112399993952099   0.592773651169898   0.25187789584633863   0.8446695323944762   0.9563859988003603   0.3527252132931679   0.9956272584269797   0.2779688896509742   0.530965406627134   0.4650071387459417   0.29235100997383784   0.8897690875972933   0.29500197181816007   0.09660506606007453
0.17865568630351975   0.9109542105111742   0.7922251297236166   0.8250066903274322   0.22691817981195367   0.3508996801979384   0.4396191548451706   0.8660387141478431   0.4632246487530966   0.5544381689430118   0.7283791554499608   0.27326506297794506   0.211346752906758   0.7097686365485357   0.7719931566496004   0.9205398496847772   0.2157194944797783   0.4317997468975615   0.24102775002246654   0.45553271093883546   0.9233684845059404   0.5420306593002682   0.9460257782043064   0.35892764487876094   0.7447127982024208   0.631076448789094   0.15380064848068992   0.5339209545513287   0.517794618390467   0.28017676859115564   0.7141814936355193   0.6678822404034855   0.054569969637370465   0.7257385996481438   0.9858023381855585   0.3946171774255405   0.8432232167306124   0.015969963099608086   0.21380918153595804   0.47407732774076333   0.6275037222508342   0.5841702162020466   0.9727814315134915   0.01854461680192786   0.7041352377448936   0.042139556901778445   0.026755653309185015   0.6596169719231669   0.9594224395424729   0.4110631081126844   0.8729550048284951   0.12569601737183825   0.44162782115200583   0.1308863395215288   0.1587735111929758   0.4578137769683527   0.3870578515146354   0.405147739873385   0.1729711730074173   0.06319659954281219   0.5438346347840229   0.3891777767737769   0.9591619914714593   0.5891192718020488
0.9163309125331888   0.8050075605717303   0.9863805599579678   0.570574655000121   0.21219567478829512   0.7628680036699519   0.9596249066487827   0.910957683076954   0.2527732352458222   0.3518048955572674   0.08666990182028766   0.7852616657051158   0.8111454140938164   0.22091855603573862   0.9278963906273119   0.3274478887367631   0.424087562579181   0.8157708161623536   0.7549252176198946   0.26425128919395097   0.8802529277951581   0.42659303938857673   0.7957632261484353   0.6751320173919021   0.9639220152619693   0.6215854788168464   0.8093826661904675   0.10455736239178112   0.7517263404736741   0.8587174751468946   0.8497577595416848   0.19359967931482705   0.49895310522785197   0.5069125795896271   0.7630878577213971   0.4083380136097112   0.6878076911340356   0.2859940235538885   0.8351914670940852   0.08089012487294811   0.2637201285548546   0.47022320739153484   0.08026624947419067   0.8166388356789972   0.38346720075969654   0.043630168002958145   0.2845030233257554   0.14150681828709505   0.41954518549772724   0.42204468918611177   0.47512035713528783   0.036949455895313926   0.6678188450240531   0.5633272140392173   0.6253625975936031   0.8433497765804868   0.16886573979620106   0.05641463444959011   0.8622747398722059   0.43501176297077565   0.48105804866216545   0.7704206108957016   0.027083272778120747   0.35412163809782754
0.21733792010731082   0.3001974035041668   0.94681702330393   0.5374828024188304   0.8338707193476143   0.25656723550120863   0.6623139999781748   0.39597598413173535   0.4143255338498871   0.8345225463150969   0.18719364284288686   0.3590265282364214   0.746506688825834   0.27119533227587966   0.5618310452492837   0.5156767516559345   0.577640949029633   0.21478069782628956   0.6995563053770778   0.0806649886851589   0.09658290036746754   0.4443600869305879   0.6724730325989571   0.7265433505873313   0.8792449802601567   0.14416268342642116   0.7256560092950269   0.18906054816850099   0.04537426091254242   0.8875954479252125   0.06334200931685227   0.7930845640367656   0.6310487270626554   0.053072901610115644   0.8761483664739654   0.43405803580034424   0.8845420382368213   0.781877569334236   0.31431732122468165   0.9183812841444098   0.30690108920718834   0.5670968715079464   0.6147610158476039   0.8377162954592509   0.21031818883972078   0.12273678457735851   0.9422879832486468   0.11117294487191948   0.33107320857956407   0.9785741011509373   0.21663197395361983   0.9221123967034185   0.28569894766702164   0.09097865322572483   0.15328996463676758   0.12902783266665285   0.6546502206043663   0.03790575161560919   0.27714159816280215   0.6949697968663086   0.770108182367545   0.2560281822813732   0.9628242769381206   0.7765885127218989
0.46320709316035663   0.6889313107734267   0.34806326109051666   0.938872217262648   0.2528889043206359   0.5661945261960682   0.40577527784186984   0.8276992723907285   0.9218156957410718   0.5876204250451309   0.18914330388825001   0.90558687568731   0.6361167480740502   0.4966417718194061   0.03585333925148243   0.7765590430206571   0.9814665274696839   0.4587360202037969   0.7587117410886802   0.08158924615434861   0.21135834510213894   0.2027078379224237   0.7958874641505598   0.30500073343244977   0.7481512519417823   0.5137765271489969   0.4478242030600431   0.36612851616980174   0.4952623476211464   0.9475820009529287   0.04204892521817326   0.5384292437790732   0.5734466518800746   0.3599615759077977   0.8529056213299232   0.6328423680917632   0.9373299038060243   0.8633198040883916   0.8170522820784408   0.856283325071106   0.9558633763363404   0.4045837838845947   0.05834054098976055   0.7746940789167575   0.7445050312342015   0.201875945962171   0.26245307683920077   0.46969334548430763   0.9963537792924192   0.688099418813174   0.8146288737791577   0.1035648293145059   0.5010914316712728   0.7405174178602455   0.7725799485609844   0.5651355855354326   0.9276447797911982   0.38055584195244774   0.9196743272310611   0.9322932174436694   0.9903148759851739   0.5172360378640561   0.10262204515262033   0.07600989237256345
0.03445149964883343   0.11265225397946141   0.04428150416285979   0.30131581345580605   0.28994646841463195   0.9107763080172904   0.781828427323659   0.8316224679714984   0.29359268912221276   0.22267688920411632   0.9671995535445014   0.7280576386569925   0.79250125745094   0.4821594713438709   0.1946196049835169   0.1629220531215598   0.8648564776597417   0.10160362939142313   0.27494527775245575   0.23062883567789033   0.8745416016745678   0.5843675915273671   0.17232323259983542   0.15461894330532688   0.8400901020257344   0.4717153375479056   0.12804172843697564   0.8533031298495208   0.5501436336111025   0.5609390295306153   0.34621330111331666   0.021680661878022495   0.25655094448888976   0.3382621403264989   0.3790137475688153   0.29362302322103   0.4640496870379498   0.856102668982628   0.18439414258529838   0.13070097009947024   0.5991932093782081   0.7544990395912049   0.9094488648328426   0.9000721344215799   0.7246516077036401   0.1701314480638379   0.7371256322330072   0.745453191116253   0.8845615056779057   0.6984161105159323   0.6090839037960315   0.8921500612667321   0.3344178720668032   0.13747708098531708   0.2628706026827149   0.8704693993887096   0.0778669275779134   0.7992149406588183   0.8838568551138996   0.5768463761676796   0.6138172405399636   0.9431122716761902   0.6994627125286013   0.4461454060682094
0.014624031161755572   0.1886132320849853   0.7900138476957586   0.5460732716466294   0.2899724234581154   0.0184817840211474   0.052888215462751395   0.8006200805303765   0.40541091778020977   0.3200656735052151   0.44380431166671985   0.9084700192636443   0.0709930457134066   0.182588592519898   0.18093370898400496   0.038000619874934694   0.9931261181354932   0.3833736518610798   0.29707685387010535   0.4611542437072551   0.3793088775955296   0.44026138018488964   0.5976141413415041   0.015008837639045695   0.364684846433774   0.2516481480999043   0.8076002936457456   0.4689355659924162   0.0747124229756586   0.23316636407875693   0.7547120781829941   0.6683154854620398   0.6693015051954488   0.9131006905735418   0.3109077665162743   0.7598454661983954   0.5983084594820423   0.7305120980536438   0.12997405753226934   0.7218448463234607   0.605182341346549   0.347138446192564   0.832897203662164   0.26069060261620564   0.22587346375101944   0.9068770660076744   0.23528306232065987   0.2456817649771599   0.8611886173172454   0.65522891790777   0.42768276867491434   0.7767461989847437   0.7864761943415868   0.4220625538290131   0.6729706904919202   0.10843071352270398   0.11717468914613799   0.5089618632554713   0.3620629239756459   0.34858524732430857   0.5188662296640958   0.7784497652018275   0.2320888664433765   0.6267404010008479
0.9136838883175467   0.4313113190092635   0.3991916627812125   0.3660497983846423   0.6878104245665273   0.5244342530015891   0.16390860046055264   0.12036803340748237   0.8266218072492818   0.869205335093819   0.7362258317856383   0.34362183442273864   0.04014561290769501   0.447142781264806   0.06325514129371815   0.2351911209000347   0.922970923761557   0.9381809180093347   0.7011922173180724   0.8866058735757261   0.40410469409746125   0.15973115280750724   0.4691033508746958   0.2598654725748782   0.4904208057799146   0.7284198337982437   0.0699116880934833   0.8938156741902359   0.8026103812133873   0.20398558079665463   0.9060030876329307   0.7734476407827535   0.9759885739641054   0.33478024570283554   0.16977725584729236   0.4298258063600149   0.9358429610564105   0.8876374644380296   0.1065221145535742   0.1946346854599802   0.012872037294853445   0.9494565464286948   0.4053298972355019   0.30802881188425413   0.6087673431973921   0.7897253936211877   0.9362265463608062   0.04816333930937591   0.1183465374174776   0.061305559822943875   0.8663148582673228   0.15434766511914003   0.3157361562040903   0.8573199790262892   0.9603117706343921   0.3809000243363865   0.3397475822399848   0.5225397333234537   0.7905345147870998   0.9510742179763716   0.40390462118357434   0.6349022688854241   0.6840124002335256   0.7564395325163914
0.3910325838887209   0.6854457224567293   0.27868250299802366   0.4484107206321373   0.7822652406913287   0.8957203288355416   0.34245595663721756   0.4002473813227614   0.6639187032738512   0.8344147690125977   0.47614109836989477   0.2458997162036214   0.3481825470697608   0.9770947899863085   0.5158293277355026   0.8649996918672349   0.008434964829776027   0.45455505666285484   0.7252948129484028   0.9139254738908633   0.6045303436462017   0.8196527877774308   0.04128241271487727   0.15748594137447186   0.21349775975748078   0.13420706532070148   0.7625999097168537   0.7090752207423345   0.431232519066152   0.23848673648515983   0.42014395307963603   0.30882783941957315   0.7673138157923008   0.4040719674725621   0.9440028547097413   0.06292812321595175   0.41913126872254003   0.4269771774862536   0.42817352697423866   0.19792843134871685   0.410696303892764   0.9724221208233987   0.7028787140258358   0.28400295745785353   0.8061659602465624   0.15276933304596801   0.6615963013109586   0.1265170160833817   0.5926682004890815   0.01856226772526653   0.8989963915941049   0.41744179534104714   0.16143568142292955   0.7800755312401066   0.4788524385144689   0.108613955921474   0.3941218656306287   0.3760035637675446   0.5348495838047276   0.04568583270552226   0.9749905969080886   0.949026386281291   0.10667605683048893   0.8477574013568054
0.5642942930153245   0.9766042654578923   0.40379734280465307   0.5637544438989519   0.7581283327687622   0.8238349324119243   0.7422010414936945   0.4372374278155702   0.16546013227968065   0.8052726646866578   0.8432046498995895   0.019795632474523032   0.004024450856751097   0.025197133446551077   0.36435221138512064   0.911181676553049   0.6099025852261224   0.6491935696790064   0.8295026275803931   0.8654958438475268   0.6349119883180339   0.7001671833977154   0.7228265707499041   0.017738442490721353   0.07061769530270927   0.7235629179398232   0.319029227945251   0.45398399859176947   0.31248936253394705   0.8997279855278989   0.5768281864515564   0.016746570776199312   0.1470292302542664   0.0944553208412411   0.7336235365519669   0.9969509383016762   0.1430047793975153   0.06925818739469002   0.3692713251668463   0.08576926174862726   0.5331021941713928   0.42006461771568354   0.5397686975864533   0.22027341790110047   0.898190205853359   0.719897434317968   0.8169421268365492   0.20253497541037913   0.8275725105506497   0.996334516378145   0.49791289889129825   0.7485509768186096   0.5150831480167027   0.09660653085024606   0.9210847124397418   0.7318044060424104   0.3680539177624363   0.002151210009004971   0.18746117588777483   0.734853467740734   0.22504913836492102   0.932893022614315   0.8181898507209285   0.6490842059921068
0.6919469441935282   0.5128284048986315   0.27842115313447524   0.4288107880910063   0.7937567383401691   0.7929309705806633   0.46147902629792603   0.2262758126806272   0.9661842277895194   0.7965964542025183   0.9635661274066277   0.4777248358620175   0.4511010797728167   0.6999899233522723   0.04248141496688602   0.7459204298196073   0.08304716201038038   0.6978387133432674   0.8550202390791112   0.011066962078873175   0.8579980236454594   0.7649456907289524   0.03683038835818266   0.3619827560867664   0.16605107945193123   0.252117285830321   0.7584092352237074   0.9331719679957601   0.3722943411117621   0.45918631524965764   0.2969302089257814   0.706896155315133   0.40611011332224267   0.6625898610471392   0.33336408151915364   0.22917131945311534   0.955009033549426   0.962599937694867   0.29088266655226763   0.48325088963350815   0.8719618715390456   0.2647612243515996   0.43586242747315646   0.47218392755463495   0.013963847893586224   0.4998155336226472   0.39903203911497376   0.11020117146786858   0.847912768441655   0.2476982477923262   0.6406228038912664   0.1770292034721085   0.4756184273298929   0.7885119325426685   0.34369259496548493   0.4701330481569756   0.0695083140076502   0.12592207149552925   0.010328513446331272   0.24096172870386026   0.1144992804582242   0.1633221338006623   0.7194458468940637   0.7577108390703521
0.2425374089191786   0.8985609094490628   0.2835834194209072   0.2855269115157172   0.22857356102559237   0.39874537582641556   0.8845513803059334   0.1753257400478486   0.38066079258393737   0.15104712803408937   0.24392857641466706   0.9982965365757401   0.9050423652540445   0.3625351954914209   0.9002359814491822   0.5281634884187645   0.8355340512463942   0.23661312399589163   0.8899074680028508   0.28720175971490425   0.72103477078817   0.07329099019522932   0.1704616211087872   0.5294909206445522   0.4784973618689915   0.1747300807461666   0.88687820168788   0.24396400912883492   0.2499238008433991   0.775984704919751   0.002326821381946626   0.06863826908098633   0.8692630082594617   0.6249375768856616   0.7583982449672796   0.07034173250524622   0.9642206430054172   0.26240238139424077   0.8581622635180974   0.5421782440864817   0.12868659175902294   0.02578925739834916   0.9682547955152466   0.2549764843715775   0.4076518209708529   0.9524982672031198   0.7977931744064594   0.7254855637270253   0.9291544591018615   0.7777681864569532   0.9109149727185794   0.48152155459819046   0.6792306582584623   0.0017834815372021941   0.9085881513366327   0.4128832855172041   0.8099676499990006   0.37684590465154055   0.15018990636935314   0.3425415530119579   0.8457470069935834   0.11444352325729974   0.2920276428512557   0.8003633089254761
0.7170604152345604   0.08865426585895059   0.3237728473360091   0.5453868245538986   0.30940859426370754   0.13615599865583075   0.5259796729295497   0.8199012608268733   0.38025413516184614   0.3583878121988775   0.6150647002109704   0.33837970622868285   0.7010234769033838   0.35660433066167535   0.7064765488743378   0.9254964207114788   0.8910558269043832   0.9797584260101347   0.5562866425049846   0.5829548676995209   0.04530881991079984   0.8653149027528351   0.2642589996537289   0.7825915587740447   0.32824840467623945   0.7766606368938844   0.9404861523177198   0.23720473422014607   0.018839810412531896   0.6405046382380537   0.41450647938817003   0.4173034733932728   0.6385856752506858   0.2821168260391762   0.7994417791771996   0.0789237671645899   0.9375621983473019   0.9255124953775008   0.0929652303028619   0.15342734645311115   0.04650637144291876   0.9457540693673661   0.5366785877978774   0.5704724787535903   0.0011975515321189243   0.08043916661453102   0.2724195881441484   0.7878809199795456   0.6729491468558795   0.30377852972064656   0.3319334358264286   0.5506761857593995   0.6541093364433476   0.6632738914825929   0.9174269564382586   0.13337271236612672   0.015523661192661822   0.38115706544341665   0.11798517726105896   0.05444894520153682   0.07796146284535985   0.45564457006591585   0.025019946958197068   0.9010215987484257
0.031455091402441085   0.5098905006985498   0.4883413591603198   0.3305491199948354   0.030257539870322158   0.42945133408401875   0.21592177101617135   0.5426682000152898   0.35730839301444267   0.1256728043633722   0.8839883351897427   0.9919920142558903   0.703199056571095   0.46239891288077933   0.9665613787514842   0.8586193018897637   0.6876753953784333   0.08124184743736264   0.8485762014904252   0.8041703566882268   0.6097139325330734   0.6255972773714468   0.8235562545322281   0.9031487579398011   0.5782588411306323   0.11570677667289705   0.33521489537190835   0.5725996379449657   0.5480013012603101   0.6862554425888783   0.11929312435573701   0.02993143792967591   0.1906929082458675   0.5605826382255061   0.23530478916599426   0.03793942367378557   0.48749385167477244   0.0981837253447268   0.2687434104145101   0.17932012178402196   0.7998184562963392   0.016941877907364157   0.42016720892408493   0.3751497650957952   0.19010452376326578   0.39134460053591735   0.5966109543918567   0.472001007155994   0.6118456826326335   0.27563782386302027   0.26139605901994845   0.8994013692110283   0.06384438137232333   0.589382381274142   0.14210293466421142   0.8694699312813524   0.8731514731264558   0.02879974304863587   0.9067981454982171   0.8315305076075669   0.3856576214516834   0.9306160177039091   0.638054735083707   0.6522103858235448
0.5858391651553442   0.9136741397965449   0.21788752615962212   0.2770606207277497   0.3957346413920784   0.5223295392606275   0.6212765717677653   0.8050596135717556   0.783888958759445   0.2466917153976073   0.3598805127478169   0.9056582443607273   0.7200445773871216   0.6573093341234653   0.21777757808360548   0.036188313079374944   0.8468931042606658   0.6285095910748294   0.31097943258538835   0.20465780547180812   0.46123548280898236   0.6978935733709204   0.6729246975016813   0.5524474196482633   0.8753963176536381   0.7842194335743754   0.4550371713420592   0.27538679892051354   0.4796616762615597   0.2618898943137479   0.8337605995742938   0.47032718534875795   0.6957727175021148   0.015198178916140576   0.4738800868264769   0.5646689409880306   0.9757281401149931   0.3578888447926753   0.25610250874287144   0.5284806279086557   0.12883503585432732   0.7293792537178458   0.9451230761574831   0.3238228224368475   0.6675995530453449   0.03148568034692552   0.2721983786558018   0.7713754027885843   0.7922032353917068   0.24726624677255007   0.8171612073137426   0.4959886038680707   0.3125415591301471   0.9853763524588022   0.9834006077394488   0.02566141851931279   0.6167688416280324   0.9701781735426617   0.5095205209129718   0.4609924775312822   0.6410407015130392   0.6122893287499863   0.25341801217010046   0.9325118496226266
0.5122056656587118   0.8829100750321405   0.30829493601261737   0.608689027185779   0.8446061126133669   0.851424394685215   0.036096557356815544   0.8373136243971948   0.05240287722166013   0.6041581479126649   0.2189353500430729   0.34132502052912406   0.739861318091513   0.6187817954538627   0.23553474230362412   0.31566360200981125   0.1230924764634807   0.648603621911201   0.7260142213906522   0.8546711244785291   0.4820517749504415   0.03631429316121466   0.4725962092205518   0.9221592748559025   0.9698461092917297   0.15340421812907415   0.16430127320793445   0.31347024767012344   0.1252399966783627   0.30197982344385915   0.1282047158511189   0.4761566232729287   0.07283711945670256   0.6978216755311942   0.909269365808046   0.13483160274380465   0.3329758013651895   0.0790398800773316   0.6737346235044219   0.8191680007339934   0.2098833249017088   0.43043625816613057   0.9477204021137696   0.9644968762554643   0.7278315499512673   0.3941219650049159   0.47512419289321783   0.04233760139956182   0.7579854406595377   0.24071774687584177   0.3108229196852834   0.7288673537294383   0.632745443981175   0.9387379234319826   0.18261820383416455   0.25271073045650966   0.5599083245244725   0.2409162479007883   0.27334883802611853   0.117879127712705   0.22693252315928297   0.1618763678234567   0.5996142145216967   0.29871112697871166
0.017049198257574154   0.7314401096573261   0.6518938124079271   0.33421425072324734   0.28921764830630686   0.33731814465241017   0.17676961951470918   0.2918766493236855   0.5312322076467692   0.09660039777656843   0.8659466998294257   0.5630092955942472   0.8984867636655941   0.15786247434458583   0.6833284959952612   0.3102985651377375   0.3385784391411216   0.9169462264437975   0.40997965796914265   0.19241943742503248   0.11164591598183866   0.7550698586203408   0.810365443447446   0.8937083104463208   0.0945967177242645   0.023629748963014684   0.15847163103951892   0.5594940597230735   0.8053790694179577   0.6863116043106045   0.9817020115248097   0.267617410399388   0.2741468617711885   0.5897112065340361   0.11575531169538399   0.7046081148051409   0.3756600981055944   0.43184873218945025   0.43242681570012276   0.3943095496674034   0.03708165896447281   0.5149025057456527   0.022447157730980095   0.20189011224237088   0.9254357429826341   0.759832647125312   0.21208171428353412   0.30818180179605004   0.8308390252583696   0.7362028981622972   0.05361008324401519   0.7486877420729765   0.025459955840411965   0.04989129385169274   0.07190807171920545   0.4810703316735885   0.7513130940692234   0.4601800873176567   0.9561527600238214   0.7764622168684476   0.375652995963629   0.02833135512820644   0.5237259443236987   0.3821526672010442
0.3385713369991562   0.5134288493825537   0.5012787865927186   0.18026255495867333   0.41313559401652206   0.7535962022572418   0.2891970723091845   0.8720807531626233   0.5822965687581524   0.017393304094944592   0.2355869890651693   0.12339301108964681   0.5568366129177404   0.9675020102432519   0.16367891734596385   0.6423226794160584   0.805523518848517   0.5073219229255952   0.20752615732214238   0.8658604625476107   0.42987052288488803   0.47899056779738874   0.6838002129984436   0.48370779534656655   0.09129918588573184   0.965561718414835   0.18252142640572502   0.3034452403878932   0.6781635918692098   0.21196551615759318   0.8933243540965405   0.43136448722526993   0.09586702311105741   0.1945722120626486   0.6577373650313713   0.30797147613562315   0.539030410193317   0.22707020181939674   0.49405844768540735   0.6656487967195648   0.7335068913448   0.7197482788938016   0.286532290363265   0.799788334171954   0.30363636845991193   0.24075771109641284   0.6027320773648214   0.31608053882538745   0.2123371825741801   0.2751959926815778   0.4202106509590963   0.012635298437494225   0.5341735907049703   0.06323047652398463   0.5268862968625557   0.5812708112122243   0.4383065675939129   0.868658264461336   0.8691489318311846   0.27329933507660115   0.8992761574005959   0.6415880626419392   0.37509048414577717   0.6076505383570364
0.16576926605579595   0.9218397837481377   0.08855819378251216   0.8078622041850824   0.862132897595884   0.6810820726517248   0.4858261164176908   0.4917816653596949   0.6497957150217039   0.40588607997014703   0.06561546545859452   0.4791463669222007   0.1156221243167336   0.3426556034461624   0.5387291685960388   0.8978755557099765   0.6773155567228207   0.4739973389848264   0.6695802367648542   0.6245762206333753   0.7780393993222249   0.8324092763428871   0.29448975261907706   0.01692568227633885   0.6122701332664289   0.9105694925947494   0.2059315588365649   0.20906347809125644   0.7501372356705449   0.22948741994302455   0.7201054424188741   0.7172818127315616   0.100341520648841   0.8236013399728775   0.6544899769602796   0.2381354458093608   0.9847193963321074   0.4809457365267151   0.11576080836424077   0.3402598900993844   0.30740383960928663   0.0069483975418886705   0.44618057159938657   0.7156836694660091   0.5293644402870619   0.17453912119900156   0.1516908189803095   0.6987579871896703   0.917094307020633   0.2639696286042521   0.9457592601437446   0.48969450909841383   0.16695707135008805   0.03448220866122759   0.22565381772487056   0.7724126963668523   0.06661555070124706   0.2108808686883501   0.571163840764591   0.5342772505574915   0.08189615436913966   0.7299351321616351   0.45540303240035024   0.19401736045810714
0.774492314759853   0.7229867346197464   0.009222460800963686   0.478333690992098   0.2451278744727912   0.5484476134207448   0.8575316418206542   0.7795757038024277   0.3280335674521582   0.28447798481649267   0.9117723816769095   0.2898811947040139   0.1610764961020702   0.24999577615526508   0.6861185639520391   0.5174684983371616   0.09446094540082316   0.03911490746691499   0.11495472318744801   0.98319124777967   0.012564791031683483   0.30917977530527996   0.6595516907870977   0.7891738873215629   0.23807247627183048   0.5861930406855336   0.6503292299861341   0.31084019632946497   0.9929446017990393   0.0377454272647888   0.7927975881654798   0.5312644925270372   0.664911034346881   0.7532674424482961   0.8810252064885703   0.24138329782302334   0.5038345382448108   0.503271666293031   0.19490664253653128   0.7239147994858618   0.40937359284398767   0.464156758826116   0.07995191934908329   0.7407235517061916   0.39680880181230416   0.15497698352083608   0.4204002285619855   0.9515496643846287   0.1587363255404737   0.5687839428353024   0.7700709985758515   0.6407094680551637   0.16579172374143444   0.5310385155705136   0.9772734104103715   0.10944497552812651   0.5008806893945534   0.7777710731222176   0.09624820392180122   0.8680616777051032   0.9970461511497426   0.2744994068291865   0.9013415613852699   0.14414687821924144
0.5876725583057549   0.8103426480030704   0.8213896420361867   0.4034233265130498   0.19086375649345075   0.6553656644822344   0.40098941347420114   0.45187366212842106   0.03212743095297702   0.08658172164693194   0.6309184148983497   0.8111641940732573   0.8663357072115426   0.5555432060764183   0.6536450044879781   0.7017192185451309   0.3654550178169892   0.7777721329542007   0.5573968005661769   0.8336575408400276   0.3684088666672466   0.5032727261250142   0.656055239180907   0.6895106626207862   0.7807363083614917   0.6929300781219437   0.8346655971447203   0.2860873361077364   0.5898725518680409   0.03756441363970931   0.4336761836705192   0.8342136739793153   0.5577451209150639   0.9509826919927774   0.8027577687721695   0.02304947990605798   0.6914094137035213   0.3954394859163591   0.14911276428419137   0.3213302613609272   0.32595439588653213   0.6176673529621584   0.5917159637180145   0.48767272052089955   0.9575455292192856   0.11439462683714419   0.9356607245371075   0.7981620579001133   0.1768092208577939   0.42146454871520045   0.10099512739238718   0.5120747217923769   0.5869366689897529   0.38390013507549114   0.667318943721868   0.6778610478130617   0.02919154807468909   0.4329174430827138   0.8645611749496984   0.6548115679070037   0.3377821343711678   0.03747795716635469   0.7154484106655071   0.3334813065460765
0.011827738484635645   0.4198106042041963   0.12373244694749261   0.845808586025177   0.05428220926535009   0.3054159773670521   0.1880717224103851   0.04764652812506362   0.8774729884075562   0.8839514286518516   0.08707659501799793   0.5355718063326866   0.2905363194178032   0.5000512935763605   0.41975765129612996   0.8577107585196251   0.2613447713431141   0.06713385049364669   0.5551964763464314   0.20289919061262138   0.9235626369719463   0.02965589332729199   0.8397480656809244   0.8694178840665449   0.9117348984873107   0.6098452891230957   0.7160156187334318   0.02360929804136794   0.8574526892219606   0.30442931175604354   0.5279438963230467   0.9759627699163044   0.9799797008144044   0.42047788310419193   0.44086730130504875   0.4403909635836177   0.6894433813966012   0.9204265895278314   0.021109650008918797   0.5826802050639927   0.4280986100534871   0.8532927390341848   0.4659131736624873   0.37978101445137125   0.5045359730815407   0.8236368457068928   0.6261651079815629   0.5103631303848263   0.59280107459423   0.21379155658379706   0.9101494892481311   0.48675383234345837   0.7353483853722694   0.9093622448277535   0.3822055929250845   0.510791062427154   0.755368684557865   0.4888843617235616   0.9413382916200357   0.0704000988435364   0.06592530316126383   0.5684577721957301   0.920228641611117   0.4877198937795438
0.6378266931077767   0.7151650331615454   0.4543154679486296   0.10793887932817256   0.133290720026236   0.8915281874546527   0.8281503599670667   0.5975757489433462   0.540489645432006   0.6777366308708556   0.9180008707189355   0.11082191659988787   0.8051412600597365   0.768374386043102   0.535795277793851   0.6000308541727338   0.04977257550187145   0.2794900243195405   0.5944569861738154   0.5296307553291975   0.9838472723406076   0.7110322521238104   0.6742283445626984   0.041910861549653636   0.34602057923283086   0.9958672189622649   0.2199128766140688   0.933971982221481   0.2127298592065949   0.10433903150761224   0.3917625166470021   0.33639623327813484   0.672240213774589   0.42660240063675664   0.4737616459280666   0.22557431667824696   0.8670989537148525   0.6582280145936545   0.9379663681342155   0.6255434625055132   0.817326378212981   0.37873799027411403   0.34350938196040015   0.09591270717631571   0.8334791058723734   0.6677057381503038   0.6692810373977017   0.054001845626662076   0.48745852663954253   0.6718385191880388   0.44936816078363295   0.120029863405181   0.2747286674329476   0.5674994876804266   0.057605644136630815   0.7836336301270462   0.6024884536583587   0.1408970870436699   0.5838439982085643   0.5580593134487992   0.7353894999435062   0.48266907245001534   0.6458776300743487   0.9325158509432862
0.9180631217305252   0.10393108217590132   0.3023682481139486   0.8366031437669704   0.08458401585815171   0.4362253440255976   0.6330872107162469   0.7826012981403083   0.5971254892186092   0.7643868248375588   0.18371904993261387   0.6625714347351274   0.32239682178566154   0.19688733715713225   0.12611340579598307   0.8789378046080811   0.7199083681273029   0.05599025011346234   0.5422694075874188   0.3208784911592819   0.9845188681837967   0.573321177663447   0.8963917775130701   0.3883626402159958   0.06645574645327158   0.4693900954875457   0.5940235293991215   0.5517594964490254   0.9818717305951199   0.03316475146194806   0.9609363186828748   0.7691581983087171   0.3847462413765107   0.26877792662438926   0.7772172687502609   0.10658676357358979   0.06234941959084916   0.071890589467257   0.6511038629542778   0.22764895896550866   0.34244105146354625   0.01590033935379466   0.10883445536685897   0.9067704678062267   0.35792218327974956   0.44257916169034767   0.21244267785378887   0.518407827590231   0.29146643682647794   0.973189066202802   0.6184191484546673   0.9666483311412055   0.3095947062313581   0.9400243147408539   0.6574828297717925   0.19749013283248845   0.9248484648548474   0.6712463881164646   0.8802655610215316   0.09090336925889866   0.8624990452639982   0.5993557986492077   0.2291616980672539   0.86325441029339
0.5200579938004519   0.583455459295413   0.12032724270039491   0.9564839424871633   0.16213581052070242   0.14087629760506534   0.9078845648466061   0.4380761148969323   0.8706693736942245   0.16768723140226333   0.28946541639193873   0.47142778375572675   0.5610746674628664   0.2276629166614094   0.6319825866201462   0.2739376509232383   0.636226202608019   0.5564165285449447   0.7517170255986145   0.18303428166433966   0.7737271573440208   0.957060729895737   0.5225553275313606   0.31977987137094965   0.2536691635435688   0.373605270600324   0.40222808483096567   0.3632959288837864   0.09153335302286637   0.23272897299525863   0.49434351998435966   0.925219813986854   0.22086397932864194   0.0650417415929953   0.2048781035924209   0.45379203023112735   0.6597893118657756   0.8373788249315859   0.5728955169722747   0.17985437930788903   0.02356310925775659   0.2809622963866412   0.8211784913736603   0.9968200976435494   0.24983595191373584   0.3239015664909042   0.29862316384229964   0.6770402262725997   0.996166788370167   0.9502962958905802   0.896395079011334   0.3137442973888133   0.9046334353473007   0.7175673228953215   0.4020515590269743   0.3885244834019592   0.6837694560186588   0.6525255813023263   0.19717345543455342   0.9347324531708319   0.0239801441528832   0.8151467563707403   0.6242779384622787   0.7548780738629428
0.0004170348951266119   0.5341844599840991   0.8030994470886185   0.7580579762193935   0.7505810829813908   0.21028289349319493   0.5044762832463189   0.08101774994679378   0.7544142946112237   0.2599865976026147   0.6080812042349849   0.7672734525579805   0.849780859263923   0.5424192747072931   0.2060296452080106   0.3787489691560213   0.16601140324526426   0.8898936934049669   0.008856189773457163   0.44401651598518943   0.14203125909238104   0.07474693703422658   0.38457825131117845   0.6891384421222466   0.14161422419725445   0.5405624770501275   0.5814788042225599   0.9310804659028531   0.3910331412158637   0.33027958355693254   0.07700252097624113   0.8500627159560593   0.63661884660464   0.07029298595431782   0.46892131674125626   0.08278926339807881   0.786837987340717   0.5278737112470246   0.26289167153324566   0.7040402942420575   0.6208265840954527   0.6379800178420577   0.2540354817597885   0.2600237782568681   0.47879532500307165   0.5632330808078312   0.86945723044861   0.5708853361346216   0.3371811008058172   0.0226706037577037   0.2879784262260501   0.6398048702317685   0.9461479595899536   0.6923910202007711   0.21097590524980891   0.7897421542757092   0.3095291129853136   0.6220980342464534   0.7420545885085527   0.7069528908776304   0.5226911256445966   0.09422432299942869   0.479162916975307   0.002912596635572807
0.901864541549144   0.45624430515737097   0.22512743521551853   0.7428888183787047   0.42306921654607227   0.8930112243495398   0.35567020476690847   0.17200348224408318   0.08588811574025507   0.870340620591836   0.06769177854085842   0.5321986120123148   0.13974015615030153   0.17794960039106492   0.8567158732910495   0.7424564577366056   0.830211043164988   0.5558515661446116   0.11466128478249682   0.03550356685897526   0.30751991752039126   0.4616272431451829   0.6354983678071898   0.03259097022340245   0.40565537597124735   0.005382937987811951   0.4103709325916713   0.2897021518446977   0.982586159425175   0.11237171363827217   0.0547007278247628   0.11769866960061456   0.89669804368492   0.24203109304643608   0.9870089492839044   0.5855000575882998   0.7569578875346185   0.06408149265537116   0.13029307599285486   0.8430435998516942   0.9267468443696305   0.5082299265107596   0.015631791210358053   0.807540032992719   0.6192269268492393   0.04660268336557669   0.38013342340316825   0.7749490627693165   0.21357155087799193   0.04121974537776474   0.969762490811497   0.4852469109246188   0.23098539145281688   0.9288480317394926   0.9150617629867341   0.3675482413240042   0.3342873477678969   0.6868169386930565   0.9280528137028298   0.7820481837357044   0.5773294602332785   0.6227354460376853   0.7977597377099749   0.9390045838840101
0.6505826158636479   0.11450551952692573   0.7821279464996168   0.13146455089129114   0.03135568901440863   0.06790283616134904   0.4019945230964486   0.3565154881219746   0.8177841381364167   0.0266830907835843   0.43223203228495166   0.8712685771973558   0.5867987466835998   0.09783505904409173   0.5171702692982175   0.5037203358733516   0.2525113989157029   0.41101812035103524   0.5891174555953876   0.7216721521376472   0.6751819386824245   0.78828267431335   0.7913577178854128   0.782667568253637   0.024599322818776553   0.6737771547864242   0.009229771385795917   0.651203017362346   0.993243633804368   0.6058743186250751   0.6072352482893473   0.29468752924037134   0.17545949566795122   0.5791912278414909   0.17500321600439567   0.4234189520430155   0.5886607489843514   0.4813561687973991   0.6578329467061782   0.9196986161696639   0.3361493500686485   0.07033804844636388   0.06871549111079048   0.19802646403201665   0.6609674113862241   0.28205537413301396   0.2773577732253777   0.4153588957783796   0.6363680885674475   0.6082782193465898   0.2681280018395818   0.7641558784160336   0.6431244547630796   0.0024039007215145803   0.6608927535502345   0.4694683491756623   0.46766495909512834   0.42321267288002373   0.4858895375458388   0.04604939713264681   0.8790042101107769   0.9418565040826246   0.8280565908396607   0.1263507809629829
0.5428548600421285   0.8715184556362607   0.7593410997288702   0.9283243169309663   0.8818874486559044   0.5894630815032468   0.48198332650349246   0.5129654211525867   0.24551936008845687   0.981184862156657   0.2138553246639107   0.7488095427365531   0.6023949053253773   0.9787809614351425   0.5529625711136762   0.27934119356089077   0.13472994623024892   0.5555682885551187   0.06707303356783739   0.23329179642824396   0.25572573611947197   0.6137117844724941   0.23901644272817674   0.10694101546526102   0.7128708760773436   0.7421933288362335   0.4796753429993066   0.17861669853429477   0.8309834274214392   0.15273024733298665   0.9976920164958141   0.665651277381708   0.5854640673329823   0.17154538517632964   0.7838366918319034   0.916841734645155   0.9830691620076051   0.19276442374118719   0.2308741207182272   0.6375005410842642   0.8483392157773562   0.6371961351860684   0.16380108715038977   0.40420874465602025   0.5926134796578841   0.023484350713574326   0.9247846444222131   0.2972677291907592   0.8797426035805406   0.2812910218773409   0.44510930142290644   0.11865103065646448   0.04875917615910141   0.12856077454435424   0.4474172849270924   0.4529997532747564   0.4632951088261191   0.9570153893680247   0.663580593095189   0.5361580186296014   0.48022594681851405   0.7642509656268375   0.4327064723769618   0.8986574775453372
0.6318867310411579   0.12705483044076898   0.268905385226572   0.4944487328893169   0.0392732513832738   0.10357047972719466   0.34412074080435895   0.19718100369855768   0.1595306478027332   0.8222794578498538   0.8990114393814526   0.0785299730420932   0.11077147164363181   0.6937186833054995   0.45159415445436013   0.6255302197673368   0.6474763628175128   0.7367032939374749   0.7880135613591712   0.08937220113773536   0.16725041599899867   0.9724523283106374   0.3553070889822094   0.19071472359239816   0.5353636849578407   0.8453974978698685   0.0864017037556374   0.6962659907030813   0.49609043357456695   0.7418270181426738   0.7422809629512784   0.4990849870045236   0.3365597857718337   0.91954756029282   0.8432695235698259   0.42055501396243034   0.2257883141282019   0.22582887698732057   0.39167536911546574   0.7950247941950935   0.5783119513106892   0.48912558304984566   0.6036618077562945   0.7056525930573582   0.41106153531169054   0.5166732547392082   0.24835471877408516   0.51493786946496   0.8756978503538498   0.6712757568693398   0.16195301501844778   0.8186718787618787   0.37960741677928284   0.929448738726666   0.41967205206716934   0.3195868917573552   0.04304763100744913   0.009901178433845935   0.5764025284973434   0.8990318777949249   0.8172593168792472   0.7840723014465254   0.1847271593818777   0.10400708359983131
0.238947365568558   0.2949467183966797   0.5810653516255831   0.3983544905424731   0.8278858302568675   0.7782734636574714   0.332710632851498   0.8834166210775131   0.9521879799030176   0.10699770678813166   0.17075761783305018   0.06474474231563433   0.5725805631237348   0.17754896806146567   0.7510855657658808   0.7451578505582791   0.5295329321162857   0.16764778962761973   0.1746830372685374   0.8461259727633542   0.7122736152370385   0.3835754881810943   0.9899558778866597   0.742118889163523   0.47332624966848047   0.08862876978441465   0.4088905262610765   0.34376439862104985   0.645440419411613   0.31035530612694323   0.07617989340957858   0.46034777754353673   0.6932524395085954   0.20335759933881156   0.9054222755765284   0.39560303522790236   0.12067187638486052   0.025808631277345905   0.15433670981064754   0.6504451846696232   0.5911389442685748   0.8581608416497262   0.9796536725421101   0.804319211906269   0.8788653290315364   0.47458535346863184   0.9896977946554505   0.06220032274274605   0.40553907936305583   0.3859565836842172   0.5808072683943739   0.7184359241216962   0.7600986599514429   0.07560127755727396   0.5046273749847954   0.25808814657815954   0.06684622044284749   0.8722436782184624   0.5992050994082669   0.8624851113502572   0.946174344057987   0.8464350469411165   0.4448683895976194   0.2120399266806339
0.3550353997894122   0.9882742052913903   0.46521471705550926   0.4077207147743649   0.4761700707578758   0.5136888518227585   0.4755169224000588   0.34552039203161883   0.07063099139481999   0.1277322681385413   0.8947096540056848   0.6270844679099227   0.31053233144337716   0.05213099058126734   0.3900822790208895   0.36899632133176313   0.24368611100052967   0.17988731236280495   0.7908771796126226   0.506511209981506   0.29751176694254267   0.33345226542168843   0.3460087900150032   0.2944712833008721   0.9424763671531305   0.3451780601302981   0.880794072959494   0.8867505685265072   0.46630629639525467   0.8314892083075397   0.40527715055943514   0.5412301764948884   0.3956753050004347   0.7037569401689984   0.5105674965537503   0.9141457085849657   0.08514297355705754   0.651625949587731   0.12048521753286082   0.5451493872532026   0.8414568625565279   0.4717386372249261   0.32960803792023824   0.038638177271696626   0.5439450956139852   0.13828637180323763   0.9835992479052351   0.7441668939708246   0.6014687284608546   0.7931083116729395   0.10280517494574119   0.8574163254443173   0.1351624320656   0.9616191033653998   0.697528024386306   0.31618614894942904   0.7394871270651653   0.2578621631964015   0.1869605278325557   0.4020404403644633   0.6543441535081078   0.6062362136086705   0.0664753102996949   0.8568910531112607
0.8128872909515799   0.1344975763837444   0.7368672723794566   0.8182528758395641   0.26894219533759467   0.9962112045805068   0.7532680244742216   0.07408598186873952   0.66747346687674   0.2031028929075673   0.6504628495284803   0.21666965642442218   0.53231103481114   0.24148378954216745   0.9529348251421743   0.9004835074749932   0.7928239077459747   0.983621626345766   0.7659742973096186   0.4984430671105299   0.1384797542378669   0.3773854127370955   0.6994989870099237   0.6415520139992692   0.32559246328628705   0.2428878363533511   0.962631714630467   0.8232991381597051   0.056650267948692344   0.2466766317728443   0.2093636901562455   0.7492131562909656   0.38917680107195235   0.04357373886527701   0.5589008406277651   0.5325434998665435   0.8568657662608123   0.8020899493231095   0.6059660154855908   0.6320599923915503   0.06404185851483768   0.8184683229773435   0.8399917181759723   0.1336169252810204   0.9255621042769707   0.44108291024024804   0.14049273116604855   0.4920649112817512   0.5999696409906837   0.19819507388689697   0.1778610165355815   0.6687657731220461   0.5433193730419914   0.9515184421140527   0.9684973263793359   0.9195526168310805   0.15414257197003903   0.9079447032487756   0.4095964857515708   0.3870091169645371   0.29727680570922665   0.10585475392566611   0.80363047026598   0.7549491245729868
0.233234947194389   0.28738643094832256   0.9636387520900077   0.6213321992919664   0.30767284291741825   0.8463035207080745   0.8231460209239592   0.1292672880102152   0.7077032019267345   0.6481084468211775   0.6452850043883777   0.4605015148881691   0.1643838288847431   0.6965900047071248   0.6767876780090416   0.5409488980570886   0.010241256914704067   0.7886453014583492   0.26719119225747084   0.1539397810925515   0.7129644512054774   0.6827905475326831   0.4635607219914909   0.39899065651956467   0.4797295040110884   0.39540411658436053   0.4999219699014832   0.7776584572275983   0.17205666109367015   0.5491005958762861   0.676775948977524   0.648391169217383   0.46435345916693566   0.9009921490551086   0.03149094458914638   0.18788965432921395   0.2999696302821926   0.2044021443479837   0.3547032665801047   0.6469407562721253   0.2897283733674885   0.4157568428896345   0.08751207432263389   0.49300097517957386   0.5767639221620111   0.7329662953569515   0.623951352331143   0.09401031866000921   0.09703441815092272   0.33756217877259087   0.12402938242965984   0.31635186143241095   0.9249777570572525   0.7884615828963047   0.4472534334521358   0.6679606922150279   0.4606242978903169   0.8874694338411963   0.41576248886298944   0.48007103788581396   0.1606546676081243   0.6830672894932125   0.06105922228288472   0.8331302816136885
0.8709262942406358   0.267310446603578   0.9735471479602509   0.3401293064341147   0.29416237207862467   0.5343441512466266   0.3495957956291078   0.24611898777410549   0.19712795392770197   0.19678197247403575   0.22556641319944798   0.9297671263416946   0.27215019687044945   0.408320389577731   0.7783129797473122   0.26180643412666665   0.8115258989801326   0.5208509557365347   0.36255049088432273   0.7817353962408526   0.6508712313720083   0.8377836662433222   0.301491268601438   0.9486051146271641   0.7799449371313725   0.5704732196397442   0.32794412064118716   0.6084758081930495   0.48578256505274775   0.036129068393117546   0.9783483250120794   0.36235682041894396   0.28865461112504576   0.8393470959190817   0.7527819118126313   0.43258969407724945   0.01650441425459635   0.4310267063413508   0.9744689320653191   0.1707832599505828   0.20497851527446379   0.9101757506048161   0.6119184411809965   0.3890478637097301   0.5541072839024556   0.07239208436149393   0.3104271725795585   0.440442749082566   0.7741623467710831   0.5019188647217497   0.9824830519383713   0.8319669408895165   0.28837978171833534   0.4657897963286322   0.004134726926291973   0.46961012047057255   0.9997251705932896   0.6264427004095504   0.2513528151136606   0.03702042639332314   0.9832207563386932   0.1954159940681996   0.27688388304834144   0.8662371664427403
0.7782422410642295   0.28524024346338345   0.664965441867345   0.47718930273301025   0.22413495716177387   0.21284815910188953   0.3545382692877865   0.03674655365044425   0.4499726103906908   0.7109292943801397   0.37205521734941516   0.2047796127609277   0.16159282867235547   0.24513949805150756   0.3679204904231232   0.7351694922903551   0.16186765807906592   0.6186967976419572   0.11656767530946256   0.698149065897032   0.17864690174037273   0.4232808035737576   0.8396837922611211   0.8319118994542917   0.40040466067614333   0.13804056011037408   0.1747183503937762   0.3547225967212814   0.17626970351436946   0.9251924010084845   0.8201800811059897   0.3179760430708372   0.7262970931236786   0.21426310662834477   0.44812486375657457   0.11319643030990947   0.5647042644513232   0.9691236085768372   0.0802043733334514   0.37802693801955434   0.40283660637225727   0.3504268109348801   0.9636366980239889   0.6798778721225224   0.22418970463188456   0.9271460073611225   0.12395290576286769   0.8479659726682307   0.8237850439557413   0.7891054472507484   0.9492345553690915   0.4932433759469492   0.6475153404413718   0.8639130462422638   0.12905447426310176   0.17526733287611201   0.9212182473176931   0.6496499396139191   0.6809296105065272   0.06207090256620255   0.3565139828663699   0.6805263310370819   0.6007252371730758   0.6840439645466482
0.9536773764941127   0.33009952010220184   0.6370885391490869   0.004166092424125885   0.7294876718622281   0.40295351274107927   0.5131356333862193   0.15620011975589523   0.9057026279064868   0.6138480654903309   0.5639010780171277   0.662956743808946   0.25818728746511505   0.7499350192480669   0.434846603754026   0.48768941093283397   0.3369690401474219   0.10028507963414786   0.7539169932474988   0.42561850836663145   0.980455057281052   0.41975874859706597   0.15319175607442304   0.7415745438199832   0.026777680786939352   0.08965922849486414   0.5161032169253361   0.7374084513958573   0.2972900089247113   0.6867057157537848   0.0029675835391168785   0.5812083316399621   0.3915873810182245   0.072857650263454   0.4390665055219891   0.9182515878310161   0.13340009355310944   0.32292263101538704   0.004219901767963147   0.4305621768981821   0.7964310534056875   0.22263755138123917   0.25030290852046433   0.004943668531550684   0.8159759961246356   0.8028788027841732   0.09711115244604128   0.2633691247115675   0.7891983153376962   0.713219574289309   0.5810079355207052   0.5259606733157102   0.49190830641298494   0.0265138585355242   0.5780403519815883   0.9447523416757481   0.10032092539476045   0.9536562082720702   0.13897384645959915   0.026500753844731918   0.966920831841651   0.6307335772566832   0.134753944691636   0.5959385769465498
0.17048977843596347   0.408096025875444   0.8844510361711717   0.5909949084149991   0.3545137823113279   0.6052172230912708   0.7873398837251304   0.32762578370343165   0.5653154669736317   0.8919976488019618   0.20633194820442521   0.8016651103877215   0.07340716056064679   0.8654837902664375   0.6282915962228369   0.8569127687119735   0.9730862351658863   0.9118275819943673   0.4893177497632378   0.8304120148672416   0.006165403324235329   0.2810940047376842   0.35456380507160173   0.23447343792069178   0.8356756248882719   0.8729979788622402   0.4701127689004301   0.6434785295056926   0.48116184257694394   0.2677807557709694   0.6827728851752997   0.315852745802261   0.9158463756033123   0.37578310696900763   0.4764409369708745   0.5141876354145395   0.8424392150426654   0.5102993167025701   0.8481493407480375   0.657274866702566   0.8693529798767791   0.5984717347082028   0.3588315909847998   0.8268628518353244   0.8631875765525437   0.3173777299705186   0.004267785913198005   0.5923894139146326   0.02751195166427191   0.44437975110827843   0.5341550170127679   0.94891088440894   0.546350109087328   0.17659899533730902   0.8513821318374682   0.6330581386066789   0.6305037334840158   0.8008158883683014   0.3749411948665938   0.11887050319213945   0.7880645184413503   0.2905165716657313   0.5267918541185562   0.46159563648957347
0.9187115385645712   0.6920448369575285   0.16796026313375648   0.6347327846542491   0.05552396201202744   0.3746671069870099   0.16369247722055846   0.04234337073961644   0.028012010347755526   0.9302873558787315   0.6295374602077906   0.0934324863306765   0.48166190126042757   0.7536883605414225   0.7781553283703223   0.46037434772399755   0.8511581677764118   0.9528724721731211   0.40321413350372853   0.3415038445318581   0.06309364933506151   0.6623559005073898   0.8764222793851723   0.8799082080422846   0.14438211077049032   0.9703110635498613   0.7084620162514158   0.24517542338803558   0.08885814875846287   0.5956439565628514   0.5447695390308573   0.20283205264841914   0.060846138410707344   0.6653566006841198   0.9152320788230668   0.10939956631774266   0.5791842371502798   0.9116682401426974   0.13707675045274453   0.6490252185937451   0.7280260693738679   0.9587957679695763   0.733862616949016   0.307521374061887   0.6649324200388065   0.29643986746218653   0.8574403375638437   0.4276131660196023   0.5205503092683161   0.32612880391232524   0.14897832131242786   0.18243774263156676   0.43169216050985326   0.7304848473494738   0.6042087822815705   0.9796056899831476   0.37084602209914597   0.065128246665354   0.6889767034585036   0.870206123665405   0.7916617849488662   0.15346000652265657   0.5518999530057591   0.22118090507165986
0.06363571557499818   0.19466423855308024   0.8180373360567431   0.9136595310097728   0.3987032955361917   0.8982243710908937   0.9605969984928994   0.4860463649901705   0.8781529862678756   0.5720955671785685   0.8116186771804715   0.3036086223586038   0.4464608257580223   0.8416107198290946   0.20740989489890108   0.3240029323754562   0.07561480365887636   0.7764824731637406   0.5184331914403975   0.45379680871005124   0.2839530187100102   0.6230224666410841   0.9665332384346383   0.23261590363839138   0.22031730313501202   0.4283582280880038   0.14849590237789523   0.31895637262861853   0.8216140075988203   0.5301338569971101   0.18789890388499583   0.832910007638448   0.9434610213309447   0.9580382898185416   0.37628022670452427   0.5293013852798442   0.4970001955729224   0.116427569989447   0.16887033180562316   0.20529845290438803   0.42138539191404606   0.3399450968257064   0.6504371403652257   0.7515016441943368   0.13743237320403584   0.7169226301846223   0.6839039019305874   0.5188857405559454   0.9171150700690238   0.2885644020966186   0.5354079995526921   0.19992936792732688   0.09550106247020353   0.7584305450995085   0.34750909566769633   0.3670193602888789   0.1520400411392588   0.8003922552809669   0.9712288689631721   0.8377179750090347   0.6550398455663364   0.6839646852915199   0.8023585371575489   0.6324195221046467
0.23365445365229037   0.3440195884658135   0.15192139679232317   0.8809178779103098   0.09622208044825452   0.6270969582811912   0.46801749486173577   0.36203213735436446   0.1791070103792307   0.33853255618457256   0.9326094953090436   0.16210276942703755   0.08360594790902719   0.5801020110850641   0.5851003996413473   0.7950834091381587   0.9315659067697684   0.7797097558040972   0.6138715306781752   0.957365434129124   0.276526061203432   0.09574507051257727   0.8115129935206263   0.32494591202447737   0.042871607551141604   0.7517254820467638   0.6595915967283033   0.4440280341141675   0.9466495271028871   0.12462852376557268   0.19157410186656743   0.0819958967598031   0.7675425167236564   0.7860959675810002   0.2589646065575238   0.9198931273327655   0.6839365688146292   0.2059939564959361   0.6738642069161765   0.12480971819460686   0.7523706620448608   0.426284200691839   0.05999267623800126   0.16744428406548287   0.4758446008414288   0.3305391301792617   0.2484796827173749   0.8424983720410055   0.4329729932902872   0.5788136481324979   0.5888880859890717   0.39847033792683795   0.48632346618740013   0.4541851243669252   0.39731398412250424   0.3164744411670349   0.7187809494637438   0.6680891567859251   0.13834937756498042   0.39658131383426937   0.0348443806491146   0.46209520028998896   0.4644851706488039   0.27177159563966247
0.2824737186042538   0.035810999598149984   0.40449249441080265   0.10432731157417963   0.806629117762825   0.7052718694188883   0.15601281169342776   0.26182893953317415   0.3736561244725377   0.12645822128639045   0.5671247257043561   0.8633586016063362   0.8873326582851375   0.6722730969194652   0.16981074158185183   0.5468841604393013   0.16855170882139375   0.004183940133540203   0.03146136401687141   0.15030284660503196   0.13370732817227918   0.5420887398435512   0.5669761933680675   0.8785312509653694   0.8512336095680254   0.5062777402454013   0.16248369895726483   0.7742039393911898   0.044604491805200444   0.801005870826513   0.0064708872638370545   0.5123749998580157   0.6709483673326627   0.6745476495401225   0.439346161559481   0.6490163982516796   0.7836157090475252   0.0022745526206572825   0.26953541997762914   0.10213223781237823   0.6150640002261314   0.9980906124871171   0.2380740559607577   0.9518293912073463   0.48135667205385224   0.45600187264356584   0.6710978625926902   0.07329814024197681   0.6301230624858268   0.9497241323981646   0.5086141636354254   0.299094200850787   0.5855185706806264   0.14871826157165158   0.5021432763715883   0.7867192009927713   0.9145702033479637   0.47417061203152905   0.06279711481210737   0.13770280274109173   0.1309544943004385   0.47189605941087176   0.7932616948344783   0.0355705649287135
0.5158904940743071   0.4738054469237547   0.5551876388737206   0.08374117372136722   0.03453382202045482   0.017803574280188864   0.8840897762810304   0.010443033479390403   0.40441075953462796   0.06807944188202433   0.3754756126456049   0.7113488326286034   0.8188921888540015   0.9193611803103727   0.8733323362740166   0.9246296316358321   0.9043219855060378   0.44519056827884373   0.8105352214619093   0.7869268288947404   0.7733674912055993   0.973294508867972   0.01727352662743099   0.751356263966027   0.25747699713129224   0.49948906194421727   0.46208588775371046   0.6676150902446597   0.22294317511083744   0.4816854876640284   0.5779961114726802   0.6571720567652694   0.8185324155762095   0.4136060457820041   0.20252049882707518   0.9458232241366659   0.999640226722208   0.4942448654716313   0.32918816255305855   0.02119359250083371   0.09531824121617014   0.04905429719278761   0.5186529410911493   0.23426676360609328   0.32195075001057083   0.07575978832481566   0.5013794144637184   0.4829104996400664   0.06447375287927855   0.5762707263805984   0.039293526710007895   0.8152954093954067   0.8415305777684411   0.09458523871656996   0.46129741523732776   0.15812335263013735   0.02299816219223162   0.6809791929345659   0.2587769164102526   0.2123001284934715   0.023357935470023652   0.18673432746293456   0.929588753857194   0.19110653599263777
0.9280396942538535   0.13768003027014694   0.4109358127660447   0.9568397723865445   0.6060889442432827   0.061920241945331286   0.9095563983023264   0.4739292727464781   0.5416151913640042   0.4856495155647329   0.8702628715923184   0.6586338633510714   0.7000846135955631   0.3910642768481629   0.4089654563549907   0.5005105107209341   0.6770864514033315   0.710085083913597   0.15018853994473808   0.28821038222746265   0.6537285159333078   0.5233507564506625   0.22059978608754405   0.09710384623482486   0.7256888216794543   0.38567072618051557   0.8096639733214993   0.14026407384828038   0.11959987743617156   0.32375048423518427   0.900107575019173   0.6663348011018022   0.5779846860721674   0.8381009686704514   0.02984470342685455   0.007700937750730767   0.8779000724766043   0.44703669182228845   0.6208792470718638   0.5071904270297967   0.20081362107327289   0.7369516079086914   0.4706907071271258   0.21898004480233402   0.5470851051399651   0.21360085145802885   0.25009092103958175   0.12187619856750917   0.8213962834605109   0.8279301252775133   0.4404269477180824   0.9816121247192288   0.7017964060243392   0.5041796410423289   0.5403193726989094   0.31527732361742655   0.12381171995217188   0.6660786723718776   0.5104746692720548   0.3075763858666958   0.24591164747556754   0.21904198054958915   0.8895954222001909   0.8003859588368991
0.04509802640229466   0.48209037264089777   0.41890471507306515   0.5814059140345651   0.49801292126232954   0.26848952118286895   0.16881379403348343   0.45952971546705595   0.6766166378018187   0.44055939590535564   0.7283868463154011   0.47791759074782714   0.9748202317774795   0.9363797548630267   0.1880674736164917   0.1626402671304006   0.8510085118253076   0.2703010824911491   0.6775928043444369   0.8550638812637048   0.6050968643497401   0.05125910194155991   0.787997382144246   0.05467792242680567   0.5599988379474454   0.5691687293006621   0.36909266707118077   0.47327200839224054   0.061985916685115806   0.3006792081177932   0.20027887303769737   0.013742292925184599   0.3853692788832971   0.8601198122124375   0.4718920267222963   0.5358247021773574   0.4105490471058176   0.9237400573494109   0.28382455310580457   0.37318443504695686   0.55954053528051   0.6534389748582617   0.6062317487613677   0.5181205537832521   0.95444367093077   0.6021798729167019   0.8182343666171217   0.46344263135644637   0.3944448329833246   0.03301114361603977   0.4491416995459409   0.9901706229642058   0.3324589162982088   0.7323319354982466   0.24886282650824357   0.9764283300390212   0.9470896374149117   0.872212123285809   0.7769707997859473   0.44060362786166374   0.5365405903090942   0.9484720659363982   0.4931462466801427   0.06741919281470692
0.9770000550285841   0.29503309107813636   0.886914497918775   0.5492986390314549   0.022556384097814144   0.6928532181614345   0.06868013130165328   0.08585600767500855   0.6281115511144896   0.6598420745453947   0.6195384317557123   0.09568538471080275   0.29565263481628073   0.9275101390471482   0.3706756052474688   0.11925705467178155   0.34856299740136903   0.05529801576133911   0.5937048054615215   0.6786534268101178   0.8120224070922749   0.10682594982494094   0.1005585587813788   0.6112342339954109   0.8350223520636908   0.8117928587468045   0.2136440608626038   0.061935594963955974   0.8124659679658767   0.11893964058537007   0.14496392956095053   0.9760795872889474   0.1843544168513871   0.45909756603997537   0.5254254978052382   0.8803942025781447   0.8887017820351063   0.5315874269928272   0.15474989255776941   0.7611371479063631   0.5401387846337373   0.4762894112314881   0.5610450870962479   0.08248372109624535   0.7281163775414624   0.3694634614065471   0.46048652831486914   0.4712494871008345   0.8930940254777716   0.5576706026597426   0.24684246745226532   0.4093138921368785   0.08062805751189499   0.4387309620743725   0.10187853789131479   0.4332343048479311   0.8962736406605079   0.9796333960343971   0.5764530400860766   0.5528401022697864   0.00757185862540154   0.44804596904156996   0.4217031475283072   0.7917029543634232
0.4674330739916642   0.9717565578100819   0.8606580604320593   0.709219233267178   0.7393166964502018   0.6022930964035347   0.40017153211719014   0.23796974616634342   0.8462226709724302   0.044622493743792145   0.15332906466492485   0.828655854029465   0.7655946134605353   0.6058915316694197   0.051450526773610054   0.3954215491815338   0.8693209728000273   0.6262581356350224   0.47499748668753344   0.8425814469117474   0.8617491141746257   0.1782121665934525   0.05329433915922625   0.0508784925483242   0.39431604018296157   0.2064556087833706   0.192636278727167   0.3416592592811463   0.6549993437327597   0.6041625123798359   0.7924647466099768   0.10368951311480289   0.8087766727603296   0.5595400186360437   0.639135681945052   0.27503365908533794   0.04318205929979435   0.9536484869666241   0.5876851551714419   0.8796121099038041   0.17386108649976703   0.32739035133160166   0.11268766848390846   0.037030662992056665   0.31211197232514126   0.14917818473814914   0.059393329324682206   0.9861521704437325   0.9177959321421797   0.9427225759547785   0.8667570505975152   0.6444929111625861   0.26279658840941994   0.33856006357494267   0.07429230398753842   0.5408033980477833   0.4540199156490904   0.7790200449388989   0.43515662204248645   0.2657697389624453   0.41083785634929604   0.8253715579722748   0.8474714668710446   0.3861576290586412
0.23697676984952903   0.4979812066406732   0.734783798387136   0.3491269660665845   0.9248647975243878   0.348803021902524   0.6753904690624539   0.36297479562285206   0.007068865382208078   0.40608044594774545   0.8086334184649386   0.718481884460266   0.7442722769727881   0.06752038237280282   0.7343411144774002   0.17767848641248263   0.2902523613236977   0.2885003374339039   0.2991844924349138   0.9119087474500374   0.8794145049744017   0.4631287794616291   0.4517130255638693   0.5257511183913961   0.6424377351248727   0.965147572820956   0.7169292271767331   0.1766241523248116   0.7175729376004849   0.6163445509184319   0.04153875811427931   0.8136493567019595   0.7105040722182768   0.21026410497068643   0.23290533964934065   0.09516747224169363   0.9662317952454886   0.14274372259788362   0.49856422517194043   0.917488985829211   0.6759794339217909   0.8542433851639797   0.19937973273702664   0.005580238379173681   0.7965649289473893   0.3911146057023506   0.7476667071731574   0.47982911998777755   0.15412719382251663   0.4259670328813947   0.030737479996424195   0.30320496766296595   0.4365542562220318   0.8096224819629628   0.9891987218821449   0.4895556109610064   0.726050184003755   0.5993583769922763   0.7562933822328042   0.3943881387193128   0.7598183887582663   0.45661465439439275   0.2577291570608638   0.4768991528901018
0.08383895483647541   0.6023712692304131   0.05834942432383717   0.4713189145109281   0.2872740258890861   0.2112566635280624   0.3106827171506798   0.9914897945231506   0.1331468320665695   0.7852896306466677   0.2799452371542556   0.6882848268601846   0.6965925758445377   0.975667148683705   0.2907465152721107   0.1987292158991782   0.9705423918407827   0.37630877169142857   0.5344531330393065   0.8043410771798654   0.21072400308251632   0.9196941172970359   0.27672397597844267   0.3274419242897636   0.1268850482460409   0.3173228480666228   0.2183745516546055   0.8561230097788355   0.8396110223569547   0.10606618453856038   0.9076918345039258   0.8646332152556849   0.7064641902903853   0.32077655389189264   0.6277465973496701   0.1763483883955003   0.009871614445847594   0.3451094052081877   0.3370000820775594   0.9776191724963221   0.03932922260506491   0.9688006335167592   0.802546949038253   0.17327809531645674   0.8286052195225486   0.04910651621972333   0.5258229730598102   0.8458361710266932   0.7017201712765077   0.7317836681531006   0.30744842140520473   0.9897131612478577   0.8621091489195529   0.6257174836145402   0.39975658690127897   0.12507994599217276   0.1556449586291676   0.3049409297226475   0.7720099895516088   0.9487315575966725   0.14577334418332   0.9598315245144597   0.43500990747404944   0.9711123851003504
0.1064441215782551   0.9910308909977006   0.6324629584357966   0.7978342897838936   0.2778389020557065   0.9419243747779773   0.10663998537598632   0.9519981187572004   0.5761187307791988   0.21014070662487674   0.7991915639707816   0.9622849575093427   0.7140095818596459   0.5844232230103366   0.3994349770695026   0.83720501151717   0.5583646232304783   0.2794822932876891   0.6274249875178938   0.8884734539204976   0.4125912790471583   0.3196507687732293   0.19241508004384428   0.9173610688201472   0.30614715746890325   0.3286198777755287   0.5599521216080477   0.11952677903625362   0.028308255413196728   0.3866955029975514   0.45331213623206146   0.16752866027905317   0.45218952463399786   0.17655479637267468   0.6541205722612798   0.2052437027697104   0.738179942774352   0.5921315733623381   0.25468559519177725   0.3680386912525404   0.1798153195438736   0.31264928007464904   0.6272606076738835   0.4795652373320428   0.7672240404967152   0.9929985113014198   0.4348455276300392   0.5622041685118956   0.461076883027812   0.6643786335258911   0.8748934060219915   0.44267738947564195   0.43276862761461526   0.27768313052833965   0.42158126978993   0.2751487291965888   0.9805791029806175   0.10112833415566497   0.7674606975286502   0.0699050264268784   0.24239916020626548   0.5089967607933269   0.512775102336873   0.701866335174338
0.06258384066239188   0.1963474807186778   0.8855144946629895   0.22230109784229518   0.29535980016567664   0.20334896941725802   0.4506689670329503   0.6600969293303995   0.8342829171378646   0.538970335891367   0.5757755610109588   0.2174195398547576   0.4015142895232493   0.2612872053630273   0.15419429122102882   0.9422708106581688   0.4209351865426319   0.16015887120736236   0.38673359369237864   0.8723657842312904   0.17853602633636645   0.6511621104140355   0.8739584913555056   0.1704994490569524   0.11595218567397457   0.45481462969535774   0.9884439966925161   0.9481983512146572   0.8205923855082979   0.2514656602780997   0.5377750296595659   0.28810142188425764   0.9863094683704333   0.7124953243867327   0.9619994686486071   0.07068188202950003   0.584795178847184   0.4512081190237054   0.8078051774275782   0.12841107137133123   0.16385999230455212   0.29104924781634306   0.4210715837351996   0.2560452871400408   0.9853239659681857   0.6398871374023075   0.5471130923796939   0.08554583808308841   0.8693717802942111   0.1850725077069498   0.5586690956871777   0.13734748686843118   0.04877939478591318   0.9336068474288501   0.020894066027611808   0.8492460649841735   0.06246992641547983   0.2211115230421174   0.058894597379004765   0.7785641829546736   0.4776747475682958   0.769903404018412   0.25108941995142653   0.6501531115833423
0.3138147552637437   0.47885415620206895   0.8300178362162269   0.3941078244433015   0.32849078929555797   0.8389670187997614   0.2829047438365331   0.3085619863602131   0.45911900900134683   0.6538945110928116   0.7242356481493554   0.17121449949178189   0.4103396142154337   0.7202876636639615   0.7033415821217436   0.32196843450760837   0.34786968779995386   0.49917614062184407   0.6444469847427388   0.5434042515529348   0.870194940231658   0.7292727366034321   0.3933575647913123   0.8932511399695925   0.5563801849679144   0.25041858040136317   0.5633397285750853   0.49914331552629104   0.2278893956723564   0.41145156160160173   0.2804349847385522   0.19058132916607795   0.7687703866710095   0.7575570505087902   0.5561993365891968   0.019366829674296065   0.35843077245557586   0.03726938684482871   0.8528577544674533   0.6973983951666877   0.010561084655622022   0.5380932462229846   0.20841076972471448   0.15399414361375288   0.14036614442396397   0.8088205096195525   0.8150532049334022   0.26074300364416036   0.5839859594560496   0.5584019292181894   0.2517134763583169   0.7615996881178693   0.3560965637836932   0.14695036761658764   0.9712784916197648   0.5710183589517913   0.5873261771126836   0.38939331710779745   0.41507915503056786   0.5516515292774953   0.22889540465710778   0.35212393026296873   0.5622214005631146   0.8542531341108076
0.21833432000148575   0.8140306840399841   0.35381063083840014   0.7002589904970546   0.0779681755775218   0.005210174420431564   0.538757425904998   0.43951598685289434   0.4939822161214722   0.44680824520224216   0.287043949546681   0.677916298735025   0.137885652337779   0.2998578775856545   0.3157654579269163   0.10689793978323367   0.5505594752250953   0.9104645604778571   0.9006863028963484   0.5552464105057384   0.32166407056798757   0.5583406302148883   0.33846490233323384   0.7009932763949308   0.10332975056650179   0.7443099461749042   0.9846542714948336   0.0007342858978761585   0.02536157498898   0.7390997717544726   0.4458968455898358   0.5612182990449819   0.5313793588675078   0.29229152655223045   0.15885289604315475   0.8833020003099568   0.3934937065297288   0.9924336489665759   0.8430874381162384   0.7764040605267232   0.8429342313046334   0.08196908848871887   0.94240113521989   0.22115765002098475   0.5212701607366459   0.5236284582738305   0.6039362328866562   0.5201643736260539   0.4179404101701441   0.7793185120989263   0.6192819613918226   0.5194300877281778   0.3925788351811641   0.04021874034445375   0.17338511580198676   0.9582117886831959   0.8611994763136563   0.7479272137922233   0.014532219758831988   0.0749097883732391   0.4677057697839275   0.7554935648256473   0.17144478164259352   0.29850572784651597
0.624771538479294   0.6735244763369285   0.2290436464227035   0.07734807782553123   0.10350137774264814   0.1498960180630979   0.6251074135360473   0.5571837041994773   0.6855609675725041   0.37057750596417155   0.005825452144224759   0.03775361647129957   0.2929821323913399   0.3303587656197178   0.832440336342238   0.07954182778810366   0.4317826560776836   0.5824315518274945   0.817908116583406   0.004632039414864559   0.9640768862937561   0.8269379870018472   0.6464633349408125   0.7061263115683486   0.33930534781446203   0.15341351066491865   0.417419688518109   0.6287782337428174   0.23580397007181392   0.003517492601820723   0.7923122749820617   0.07159452954334006   0.5502430024993099   0.6329399866376492   0.786486822837837   0.033840913072040485   0.25726087010797   0.3025812210179314   0.954046486495599   0.9542990852839368   0.8254782140302864   0.7201496691904369   0.13613836991219294   0.9496670458690722   0.8614013277365303   0.8932116821885898   0.48967503497138043   0.24354073430072368   0.5220959799220682   0.7397981715236711   0.07225534645327145   0.6147625005579063   0.2862920098502543   0.7362806789218505   0.2799430714712097   0.5431679710145663   0.7360490073509444   0.10334069228420123   0.49345624863337273   0.5093270579425258   0.4787881372429744   0.8007594712662698   0.5394097621377738   0.5550279726585889
0.653309923212688   0.08060980207583293   0.40327139222558084   0.6053609267895167   0.7919085954761578   0.18739811988724314   0.9135963572542004   0.361820192488793   0.26981261555408953   0.44759994836357203   0.8413410108009289   0.7470576919308867   0.9835206057038353   0.7113192694417216   0.5613979393297193   0.20388972091632043   0.24747159835289084   0.6079785771575204   0.0679416906963465   0.6945626629737947   0.7686834611099164   0.8072191058912506   0.5285319285585727   0.13953469031520577   0.11537353789722837   0.7266093038154177   0.12526053633299192   0.5341737635256891   0.3234649424210706   0.5392111839281745   0.21166417907879154   0.17235357103689614   0.05365232686698105   0.09161123556460246   0.3703231682778626   0.42529587910600947   0.07013172116314581   0.38029196612288085   0.8089252289481433   0.22140615818968903   0.8226601228102549   0.7723133889653605   0.7409835382517969   0.5268434952158944   0.053976661700338546   0.9650942830741099   0.21245160969322416   0.3873088049006886   0.9386031238031102   0.23848497925869228   0.08719107336023224   0.8531350413749995   0.6151381813820396   0.6992737953305178   0.8755268942814407   0.6807814703381033   0.5614858545150585   0.6076625597659153   0.5052037260035781   0.25548559123209386   0.49135413335191275   0.22737059364303447   0.6962784970554348   0.03407943304240483
0.6686940105416578   0.455057204677674   0.9552949588036379   0.5072359378265104   0.6147173488413192   0.4899629216035641   0.7428433491104137   0.1199271329258219   0.6761142250382091   0.25147794234487186   0.6556522757501815   0.26679209155082245   0.060976043656169446   0.552204147014354   0.7801253814687408   0.5860106212127191   0.49949018914111093   0.9445415872484387   0.2749216554651627   0.3305250299806253   0.0081360557891982   0.7171709936054043   0.5786431584097279   0.2964455969382204   0.33944204524754046   0.2621137889277303   0.62334819960609   0.7892096591117099   0.7247246964062213   0.7721508673241662   0.8805048504956763   0.669282526185888   0.048610471368012206   0.5206729249792943   0.22485257474549483   0.4024904346350656   0.9876344277118427   0.9684687779649402   0.44472719327675403   0.8164798134223465   0.48814423857073186   0.0239271907165015   0.16980553781159138   0.48595478344172127   0.4800081827815336   0.3067561971110972   0.5911623794018634   0.18950918650350085   0.1405661375339932   0.044642408183366934   0.9678141797957734   0.4002995273917909   0.41584144112777194   0.27249154085920074   0.08730932930009715   0.7310170012059028   0.3672309697597598   0.7518186158799064   0.8624567545546024   0.32852656657083723   0.379596542047917   0.7833498379149662   0.41772956127784827   0.5120467531484908
0.8914523034771852   0.7594226471984646   0.2479240234662569   0.026091969706769493   0.4114441206956515   0.45266645008736744   0.6567616440643934   0.8365827832032686   0.2708779831616583   0.40802404190400055   0.68894746426862   0.43628325581147775   0.8550365420338863   0.13553250104479977   0.6016381349685228   0.7052662546055749   0.4878055722741266   0.38371388516489335   0.7391813804139205   0.3767396880347376   0.1082090302262096   0.6003640472499272   0.32145181913607224   0.8646929348862469   0.21675672674902446   0.8409414000514625   0.07352779566981534   0.8386009651794774   0.805312606053373   0.388274949964095   0.41676615160542196   0.002018181976208744   0.5344346228917146   0.9802509080600945   0.727818687336802   0.565734926164731   0.6793980808578283   0.8447184070152947   0.12618055236827921   0.8604686715591561   0.1915925085837017   0.46100452185040136   0.38699917195435873   0.48372898352441845   0.08338347835749209   0.8606404746004742   0.06554735281828653   0.6190360486381715   0.8666267516084676   0.019699074549011746   0.9920195571484712   0.7804350834586942   0.06131414555509468   0.6314241245849167   0.5752534055430493   0.7784169014824854   0.52687952266338   0.6511732165248223   0.8474347182062473   0.21268197531775443   0.8474814418055517   0.8064548095095275   0.721254165837968   0.35221330375859833
0.65588893322185   0.34545028765912617   0.3342549938836093   0.8684843202341799   0.572505454864358   0.48480981305865195   0.26870764106532274   0.2494482715960083   0.7058787032558904   0.46511073850964024   0.27668808391685157   0.46901318813731413   0.6445645577007957   0.8336866139247234   0.7014346783738024   0.6905962866548288   0.11768503503741563   0.18251339739990122   0.8539999601675551   0.4779143113370743   0.2702035932318639   0.37605858789037366   0.1327457943295871   0.12570100757847594   0.6143146600100138   0.030608300231247467   0.7984908004459779   0.25721668734429604   0.041809205145655816   0.5457984871725955   0.529783159380655   0.007768415748287748   0.3359305018897655   0.08068774866295528   0.2530950754638035   0.5387552276109736   0.6913659441889698   0.2470011347382318   0.5516603970900011   0.8481589409561449   0.5736809091515541   0.06448773733833058   0.6976604369224461   0.3702446296190706   0.30347731591969024   0.688429149447957   0.564914642592859   0.2445436220405947   0.6891626559096764   0.6578208492167095   0.7664238421468811   0.9873269346962986   0.6473534507640206   0.11202236204411395   0.23664068276622602   0.9795585189480109   0.3114229488742552   0.03133461338115867   0.9835456073024226   0.4408032913370373   0.6200570046852855   0.7843334786429269   0.4318852102124214   0.5926443503808924
0.04637609553373128   0.7198457413045963   0.7342247732899754   0.22239972076182174   0.742898779614041   0.03141659185663939   0.16931013069711648   0.977856098721227   0.05373612370436458   0.37359574263992995   0.4028862885502354   0.9905291640249284   0.4063826729403439   0.261573380595816   0.1662456057840094   0.010970645076917498   0.09495972406608875   0.2302387672146573   0.18269999848158688   0.5701673537398803   0.47490271938080336   0.44590528857173045   0.7508147882691655   0.9775230033589878   0.4285266238470721   0.7260595472671342   0.016590014979190097   0.7551232825971661   0.685627844233031   0.6946429554104947   0.8472798842820736   0.7772671838759391   0.6318917205286665   0.3210472127705648   0.44439359573183823   0.7867380198510107   0.22550904758832252   0.05947383217474881   0.2781479899478288   0.7757673747740932   0.13054932352223375   0.8292350649600915   0.09544799146624194   0.20560002103421293   0.6556466041414304   0.3833297763883611   0.34463320319707647   0.2280770176752251   0.22711998029435834   0.6572702291212269   0.32804318821788636   0.472953735078059   0.5414921360613273   0.9626272737107322   0.48076330393581274   0.69568655120212   0.9096004155326609   0.6415800609401674   0.03636970820397454   0.9089485313511093   0.6840913679443383   0.5821062287654186   0.7582217182561457   0.1331811565770162
0.5535420444221046   0.752871163805327   0.6627737267899038   0.9275811355428033   0.8978954402806743   0.369541387416966   0.31814052359282735   0.6995041178675782   0.6707754599863158   0.7122711582957391   0.9900973353749409   0.22655038278951917   0.12928332392498854   0.7496438845850069   0.5093340314391283   0.5308638315873991   0.21968290839232765   0.10806382364483952   0.4729643232351537   0.6219153002362898   0.5355915404479893   0.525957594879421   0.714742604979008   0.48873414365927365   0.9820494960258846   0.7730864310740938   0.05196887818910417   0.5611530081164704   0.08415405574521048   0.40354504365712784   0.7338283545962768   0.8616488902488921   0.41337859575889463   0.6912738853613887   0.7437310192213359   0.635098507459373   0.2840952718339061   0.9416300007763818   0.23439698778220763   0.10423467587197383   0.06441236344157845   0.8335661771315424   0.7614326645470539   0.482319375635684   0.5288208229935891   0.30760858225212134   0.046690059568045984   0.9935852319764104   0.5467713269677045   0.5345221511780275   0.9947211813789418   0.43243222385994   0.46261727122249396   0.13097710752089967   0.26089282678266495   0.5707833336110478   0.04923867546359935   0.43970322215951096   0.5171618075613291   0.9356848261516748   0.7651434036296932   0.49807322138312915   0.2827648197791215   0.831450150279701
0.7007310401881148   0.6645070442515868   0.5213321552320676   0.34913077464401704   0.17191021719452565   0.35689846199946546   0.47464209566402155   0.3555455426676067   0.6251388902268212   0.822376310821438   0.4799209142850797   0.9231133188076667   0.16252161900432718   0.6913992033005383   0.21902808750241473   0.3523299851966188   0.11328294354072783   0.25169598114102737   0.7018662799410856   0.416645159044944   0.3481395399110346   0.7536227597578983   0.41910146016196415   0.585195008765243   0.6474084997229198   0.08911571550631138   0.8977693049298967   0.23606423412122596   0.47549828252839416   0.7322172535068459   0.42312720926587516   0.8805186914536193   0.850359392301573   0.9098409426854079   0.9432062949807954   0.9574053726459526   0.6878377732972458   0.21844173938486963   0.7241782074783807   0.6050753874493339   0.574554829756518   0.9667457582438422   0.02231192753729505   0.18843022840438983   0.22641528984548334   0.21312299848594404   0.6032104673753309   0.6032352196391468   0.5790067901225635   0.12400728297963266   0.7054411624454342   0.36717098551792093   0.10350850759416941   0.39179002947278674   0.2823139531795591   0.4866522940643016   0.2531491152925964   0.48194908678737886   0.33910765819876365   0.529246921418349   0.5653113419953506   0.2635073474025092   0.614929450720383   0.9241715339690152
0.9907565122388328   0.29676158915866696   0.5926175231830879   0.7357413055646254   0.7643412223933493   0.0836385906727229   0.989407055807757   0.13250608592547847   0.1853344322707858   0.9596313076930902   0.2839658933623228   0.7653351004075576   0.08182592467661641   0.5678412782203035   0.0016519401827637342   0.27868280634325593   0.82867680938402   0.08589219143292463   0.6625442819840001   0.7494358849249069   0.26336546738866934   0.8223848440304155   0.0476148312636171   0.8252643509558918   0.27260895514983663   0.5256232548717484   0.4549973080805292   0.0895230453912664   0.5082677327564873   0.4419846641990256   0.4655902522727721   0.9570169594657879   0.32293330048570146   0.48235335650593536   0.1816243589104493   0.1916818590582304   0.24110737580908503   0.9145120782856319   0.17997241872768557   0.9129990527149745   0.41243056642506504   0.8286198868527073   0.5174281367436855   0.16356316779006755   0.14906509903639573   0.0062350428222918124   0.4698133054800684   0.33829881683417584   0.8764561438865591   0.4806117879505433   0.014815997399539236   0.2487757714429094   0.36818841113007184   0.03862712375151776   0.5492257451267671   0.29175881197712145   0.04525511064437041   0.5562737672455824   0.3676013862163178   0.10007695291889107   0.8041477348352853   0.6417616889599506   0.18762896748863223   0.1870779002039166
0.3917171684102203   0.8131418021072433   0.6702008307449467   0.023514732413849028   0.2426520693738246   0.8069067592849515   0.20038752526487832   0.6852159155796732   0.3661959254872655   0.32629497133440816   0.1855715278653391   0.4364401441367638   0.9980075143571936   0.2876678475828904   0.636345782738572   0.14468133215964235   0.9527524037128232   0.731394080337308   0.2687443965222542   0.04460437924075127   0.14860466887753784   0.08963239137735746   0.08111542903362196   0.8575264790368347   0.7568875004673176   0.27649058927011416   0.4109145982886752   0.8340117466229856   0.5142354310934929   0.4695838299851627   0.2105270730237969   0.14879583104331245   0.14803950560622745   0.14328885865075452   0.02495554515845781   0.7123556869065486   0.1500319912490338   0.8556210110678641   0.3886097624198858   0.5676743547469063   0.19727958753621055   0.12422693073055613   0.11986536589763165   0.523069975506155   0.04867491865867271   0.03459453935319867   0.038749936864009696   0.6655434964693203   0.2917874181913552   0.7581039500830845   0.6278353385753345   0.8315317498463347   0.7775519870978622   0.28852012009792183   0.4173082655515376   0.6827359188030222   0.6295124814916349   0.14523126144716733   0.3923527203930798   0.9703802318964736   0.47948049024260103   0.2896102503793032   0.0037429579731939455   0.4027058771495673
0.2822009027063905   0.16538331964874708   0.8838775920755623   0.8796359016434123   0.23352598404771777   0.1307887802955484   0.8451276552115526   0.21409240517409195   0.9417385658563626   0.3726848302124639   0.21729231663621812   0.38256065532775724   0.16418657875850032   0.08416471011454203   0.7999840510846805   0.699824736524735   0.5346740972668654   0.9389334486673747   0.4076313306916008   0.7294445046282614   0.05519360702426445   0.6493231982880715   0.40388837271840683   0.3267386274786941   0.7729927043178739   0.4839398786393244   0.5200107806428446   0.4471027258352818   0.5394667202701562   0.353151098343776   0.6748831254312919   0.23301032066118987   0.5977281544137937   0.9804662681313121   0.4575908087950738   0.8504496653334326   0.43354157565529333   0.89630155801677   0.6576067577103932   0.15062492880869757   0.8988674783884278   0.9573681093493953   0.2499754270187925   0.42118042418043616   0.8436738713641634   0.30804491106132387   0.8460870543003857   0.09444179670174206   0.0706811670462894   0.8241050324219995   0.32607627365754116   0.6473390708664603   0.5312144467761332   0.4709539340782235   0.6511931482262492   0.4143287502052704   0.9334862923623396   0.4904876659469114   0.19360233943117544   0.5638790848718378   0.49994471670704627   0.5941861079301413   0.5359955817207822   0.4132541560631402
0.6010772383186185   0.636817998580746   0.28602015470198966   0.992073731882704   0.7574033669544551   0.3287730875194221   0.439933100401604   0.897631935180962   0.6867221999081656   0.5046680550974226   0.11385682674406283   0.2502928643145017   0.15550775313203247   0.03371412101919912   0.4626636785178136   0.8359641141092313   0.2220214607696929   0.5432264550722877   0.26906133908663815   0.2720850292373935   0.7220767440626467   0.9490403471421465   0.733065757365856   0.8588308731742533   0.1209995057440282   0.31222234856140046   0.44704560266386634   0.8667571412915493   0.36359613878957314   0.9834492610419784   0.00711250226226235   0.9691252061105874   0.6768739388814075   0.4787812059445558   0.8932556755181995   0.7188323417960857   0.521366185749375   0.4450670849253567   0.4305919970003859   0.8828682276868544   0.29934472497968206   0.9018406298530689   0.16153065791374774   0.6107831984494608   0.5772679809170355   0.9528002827109225   0.42846490054789177   0.7519523252752075   0.4562684751730073   0.640577934149522   0.9814192978840254   0.8851951839836582   0.09267233638343413   0.6571286731075436   0.974306795621763   0.9160699778730707   0.4157983975020267   0.17834746716298783   0.08105112010356354   0.197237636076985   0.8944322117526516   0.7332803822376311   0.6504591231031777   0.3143694083901306
0.5950874867729696   0.8314397523845622   0.4889284651894299   0.7035862099406698   0.017819505855934132   0.8786394696736397   0.060463564641538126   0.9516338846654623   0.5615510306829269   0.23806153552411768   0.07904426675751272   0.06643870068180423   0.46887869429949275   0.580932862416574   0.10473747113574966   0.15036872280873353   0.053080296797466085   0.4025853952535862   0.02368635103218612   0.9531310867317485   0.1586480850448144   0.669305013015955   0.3732272279290085   0.6387616783416179   0.5635605982718448   0.8378652606313929   0.8842987627395786   0.9351754684009481   0.5457410924159107   0.9592257909577532   0.8238351980980405   0.9835415837354858   0.9841900617329838   0.7211642554336355   0.7447909313405278   0.9171028830536816   0.515311367433491   0.14023139301706142   0.6400534602047782   0.766734160244948   0.462231070636025   0.7376459977634752   0.616367109172592   0.8136030735131995   0.30358298559121055   0.06834098474752015   0.24313988124358352   0.1748413951715816   0.7400223873193658   0.2304757241161273   0.35884111850400485   0.23966592677063345   0.19428129490345505   0.2712499331583742   0.5350059204059644   0.25612434303514764   0.21009123317047124   0.5500856777247387   0.7902149890654366   0.3390214599814661   0.6947798657369801   0.4098542847076773   0.15016152886065848   0.572287299736518
0.2325487951009552   0.6722082869442021   0.5337944196880665   0.7586842262233185   0.9289658095097446   0.6038673021966819   0.29065453844448297   0.583842831051737   0.18894342219037888   0.3733915780805547   0.9318134199404781   0.3441769042811035   0.9946621272869238   0.10214164492218047   0.3968074995345137   0.08805256124595584   0.7845708941164525   0.5520559671974418   0.6065925104690771   0.7490311012644898   0.08979102837947239   0.14220168248976445   0.45643098160841866   0.1767438015279717   0.8572422332785172   0.4699933955455623   0.9226365619203521   0.41805957530465315   0.9282764237687726   0.8661260933488804   0.6319820234758692   0.8342167442529163   0.7393330015783937   0.4927345152683257   0.7001686035353911   0.4900398399718127   0.7446708742914699   0.3905928703461452   0.30336110400087746   0.4019872787258569   0.9600999801750173   0.8385369031487034   0.6967685935318003   0.6529561774613671   0.8703089517955449   0.696335220658939   0.2403376119233817   0.4762123759333954   0.01306671851702775   0.2263418251133767   0.31770105000302956   0.05815280062874223   0.08479029474825517   0.36021573176449634   0.6857190265271603   0.22393605637582603   0.34545729316986146   0.8674812164961706   0.9855504229917692   0.7338962164040134   0.6007864188783916   0.47688834615002546   0.6821893189908917   0.3319089376781565
0.6406864387033743   0.638351443001322   0.9854207254590913   0.6789527602167894   0.7703774869078293   0.9420162223423829   0.7450831135357097   0.20274038428339397   0.7573107683908016   0.7156743972290063   0.4273820635326801   0.14458758365465174   0.6725204736425463   0.35545866546450994   0.7416630370055198   0.9206515272788257   0.3270631804726849   0.4879774489683393   0.7561126140137506   0.1867553108748124   0.7262767615942933   0.01108910281831383   0.07392329502285894   0.8548463731966559   0.0855903228909191   0.37273765981699186   0.08850256956376759   0.17589361297986655   0.3152128359830898   0.4307214374746089   0.34341945602805796   0.9731532286964726   0.5579020675922883   0.7150470402456026   0.9160373924953779   0.8285656450418208   0.8853815939497419   0.35958837478109273   0.1743743554898581   0.9079141177629951   0.558318413477057   0.8716109258127535   0.41826174147610745   0.7211588068881827   0.8320416518827637   0.8605218229944397   0.3443384464532485   0.8663124336915268   0.7464513289918446   0.48778416317744777   0.25583587688948095   0.6904188207116602   0.4312384930087548   0.057062725702838886   0.9124164208614229   0.7172655920151877   0.8733364254164665   0.34201568545723626   0.9963790283660451   0.8886999469733668   0.9879548314667246   0.9824273106761435   0.822004672876187   0.9807858292103717
0.4296364179896675   0.11081638486339004   0.4037429314000795   0.259627022322189   0.5975947661069038   0.2502945618689504   0.05940448494683099   0.3933145886306622   0.8511434371150592   0.7625103986915026   0.8035686080573501   0.702895767919002   0.4199049441063044   0.7054476729886637   0.8911521871959271   0.9856301759038144   0.5465685186898379   0.36343198753142747   0.8947731588298821   0.09693022893044755   0.5586136872231133   0.381004676855284   0.07276848595369505   0.11614439972007584   0.12897726923344582   0.2701882919918939   0.6690255545536156   0.8565173773978868   0.531382503126542   0.019893730122943546   0.6096210696067845   0.4632027887672246   0.6802390660114828   0.25738333143144093   0.8060524615494344   0.7603070208482227   0.2603341219051784   0.5519356584427771   0.9149002743535074   0.7746768449444082   0.7137656032153405   0.1885036709113497   0.020127115523625366   0.6777466160139607   0.15515191599222716   0.8074989940560657   0.9473586295699303   0.5616022162938848   0.02617464675878134   0.5373107020641718   0.27833307501631477   0.705084838895998   0.49479214363223933   0.5174169719412283   0.6687120054095302   0.2418820501287734   0.8145530776207566   0.2600336405097873   0.8626595438600957   0.4815750292805508   0.5542189557155781   0.7080979820670101   0.9477592695065884   0.7068981843361425
0.8404533525002377   0.5195943111556603   0.927632153982963   0.02915156832218182   0.6853014365080105   0.7120953170995947   0.9802735244130326   0.46754935202829695   0.6591267897492291   0.1747846150354229   0.7019404493967178   0.7624645131322989   0.16433464611698978   0.6573676430941947   0.033228443987187654   0.5205824630035255   0.34978156849623326   0.3973340025844074   0.17056890012709192   0.03900743372297478   0.7955626127806551   0.6892360205173973   0.22280963062050357   0.3321092493868323   0.9551092602804175   0.16964170936173686   0.29517747663754057   0.30295768106465043   0.2698078237724071   0.4575463922621422   0.3149039522245079   0.8354083290363534   0.610681034023178   0.2827617772267193   0.61296350282779   0.07294381590405453   0.44634638790618814   0.6253941341325246   0.5797350588406024   0.552361352900529   0.0965648194099549   0.22806013154811725   0.4091661587135105   0.5133539191775542   0.3010022066292998   0.53882411103072   0.1863565280930069   0.18124466979072196   0.34589294634888224   0.36918240166898314   0.8911790514554663   0.8782869887260715   0.07608512257647515   0.911636009406841   0.5762750992309584   0.042878659689718025   0.4654040885532972   0.6288742321801216   0.9633115964031684   0.9699348437856635   0.01905770064710904   0.003480098047597005   0.38357653756256604   0.4175734908851345
0.9224928812371541   0.7754199664994798   0.9744103788490556   0.9042195717075803   0.6214906746078543   0.23659585546875975   0.7880538507560487   0.7229749019168583   0.27559772825897216   0.8674134537997766   0.8968747993005823   0.8446879131907868   0.199512605682497   0.9557774443929357   0.32059970006962396   0.8018092535010688   0.7341085171291998   0.3269032122128141   0.3572881036664556   0.8318744097154053   0.7150508164820908   0.3234231141652171   0.9737115661038895   0.4143009188302708   0.7925579352449367   0.5480031476657373   0.999301187254834   0.5100813471226905   0.17106726063708225   0.31140729219697755   0.2112473364987853   0.7871064452058322   0.8954695323781101   0.4439938383972009   0.3143725371982029   0.9424185320150453   0.695956926695613   0.4882163940042652   0.993772837128579   0.1406092785139765   0.9618484095664133   0.16131318179145115   0.6364847334621234   0.30873486879857115   0.24679759308432245   0.8378900676262341   0.6627731673582338   0.8944339499683004   0.4542396578393858   0.28988691996049676   0.6634719801033998   0.38435260284560985   0.2831723972023036   0.9784796277635192   0.4522246436046145   0.5972461576397777   0.3877028648241935   0.5344857893663183   0.1378521064064116   0.6548276256247324   0.6917459381285804   0.046269395362053024   0.14407926927783263   0.5142183471107559
0.7298975285621673   0.8849562135706018   0.5075945358157092   0.20548347831218472   0.4830999354778448   0.047066145944367796   0.8448213684574755   0.3110495283438844   0.028860277638458987   0.757179225983871   0.1813493883540756   0.9266969254982745   0.7456878804361554   0.7786995982203518   0.7291247447494611   0.32945076785849686   0.35798501561196194   0.24421380885403363   0.5912726383430494   0.6746231422337645   0.6662390774833814   0.1979444134919806   0.44719336906521684   0.1604047951230086   0.9363415489212142   0.3129881999213787   0.9395988332495075   0.9549213168108239   0.45324161344336944   0.2659220539770109   0.09477746479203214   0.6438717884669395   0.42438133580491044   0.5087428279931399   0.9134280764379565   0.7171748629686651   0.678693455368755   0.730043229772788   0.18430333168849544   0.38772409511016814   0.3207084397567931   0.48582942091875436   0.593030693345446   0.7131009528764036   0.6544693622734117   0.2878850074267738   0.1458373242802291   0.5526961577533951   0.7181278133521974   0.9748968075053951   0.2062384910307215   0.5977748409425712   0.264886199908828   0.7089747535283841   0.11146102623868936   0.9539030524756317   0.8405048641039176   0.20023192553524427   0.19803294980073283   0.23672818950696664   0.16181140873516253   0.47018869576245625   0.013729618112237389   0.8490040943967985
0.8411029689783694   0.9843592748437019   0.42069892476679144   0.13590314152039482   0.1866336067049578   0.6964742674169281   0.27486160048656233   0.5832069837669998   0.4685057933527604   0.721577459911533   0.06862310945584081   0.9854321428244286   0.20361959344393238   0.01260270638314888   0.9571620832171515   0.03152909034879692   0.3631147293400148   0.8123707808479046   0.7591291334164186   0.7948009008418303   0.20130332060485226   0.3421820850854484   0.7453995153041812   0.9457968064450318   0.36020035162648284   0.3578228102417465   0.3247005905373898   0.809893664924637   0.17356674492152502   0.6613485428248185   0.04983899005082747   0.22668668115763727   0.7050609515687647   0.9397710829132854   0.9812158805949867   0.2412545383332087   0.5014413581248323   0.9271683765301365   0.0240537973778352   0.20972544798441178   0.1383266287848175   0.11479759568223191   0.26492466396141656   0.41492454714258153   0.9370233081799653   0.7726155105967836   0.5195251486572353   0.4691277406975497   0.5768229565534824   0.414792700355037   0.19482455811984556   0.6592340757729127   0.40325621163195735   0.7534441575302187   0.14498556806901808   0.43254739461527547   0.6981952600631927   0.8136730746169332   0.16376968747403142   0.19129285628206674   0.1967539019383604   0.8865046980867967   0.13971589009619623   0.981567408297655
0.05842727315354292   0.7717071024045647   0.8747912261347797   0.5666428611550735   0.1214039649735777   0.9990915918077812   0.3552660774775443   0.09751512045752371   0.5445810084200953   0.5842988914527442   0.16044151935769876   0.438281044684611   0.14132479678813792   0.8308547339225256   0.015455951288680674   0.005733650069335556   0.4431295367249452   0.017181659305592394   0.8516862638146493   0.8144407937872689   0.2463756347865848   0.13067696121879574   0.7119703737184531   0.8328733854896139   0.18794836163304188   0.358969858814231   0.8371791475836734   0.2662305243345405   0.0665443966594642   0.35987826700644976   0.48191307010612905   0.16871540387701675   0.5219633882393689   0.7755793755537056   0.3214715507484303   0.7304343591924057   0.38063859145123097   0.94472464163118   0.30601559945974965   0.7247007091230702   0.9375090547262858   0.9275429823255876   0.45432933564510036   0.9102599153358013   0.6911334199397009   0.7968660211067919   0.7423589619266474   0.07738652984618748   0.503185058306659   0.4378961622925609   0.905179814342974   0.811156005511647   0.43664066164719484   0.07801789528611112   0.42326674423684496   0.6424406016346302   0.914677273407826   0.30243851973240554   0.10179519348841465   0.9120062424422245   0.534038681956595   0.3577138781012255   0.795779594028665   0.18730553331915437
0.5965296272303092   0.4301708957756379   0.34145025838356463   0.277045617983353   0.9053962072906083   0.633304874668846   0.5990912964569173   0.1996590881371655   0.4022111489839492   0.19540871237628507   0.6939114821139433   0.38850308262551847   0.9655704873367543   0.11739081709017395   0.2706447378770983   0.7460624809908882   0.0508932139289284   0.8149522973577684   0.16884954438868366   0.8340562385486636   0.5168545319723334   0.4572384192565429   0.37306995036001867   0.6467507052295093   0.9203249047420242   0.02706752348090507   0.03161969197645402   0.3697050872461563   0.014928697451415892   0.3937626488120591   0.43252839551953676   0.1700459991089908   0.6127175484674666   0.19835393643577404   0.7386169134055935   0.7815429164834723   0.6471470611307123   0.0809631193456001   0.46797217552849524   0.03548043549258408   0.5962538472017839   0.26601082198783166   0.2991226311398116   0.2014241969439204   0.0793993152294505   0.8087724027312887   0.926052680779793   0.5546734917144112   0.15907441048742632   0.7817048792503837   0.894432988803339   0.1849684044682548   0.14414571303601043   0.3879422304383246   0.4619045932838022   0.014922405359264023   0.5314281645685438   0.18958829400255053   0.7232876798782086   0.23337948887579174   0.8842811034378315   0.10862517465695044   0.2553155043497134   0.19789905338320765
0.2880272562360476   0.8426143526691188   0.9561928732099018   0.9964748564392872   0.20862794100659704   0.03384194993783001   0.03014019243010885   0.44180136472487613   0.049553530519170726   0.25213707068744634   0.1357072036267699   0.25683296025662133   0.9054078174831603   0.8641948402491217   0.6738026103429677   0.2419105548973573   0.37397965291461654   0.6746065462465712   0.9505149304647591   0.008531066021565559   0.4896985494767851   0.5659813715896208   0.6951994261150457   0.8106320126383579   0.20167129324073751   0.723367018920502   0.7390065529051439   0.8141571561990707   0.9930433522341404   0.689525068982672   0.708866360475035   0.37235579147419456   0.9434898217149698   0.4373879982952257   0.5731591568482651   0.11552283121757324   0.03808200423180944   0.5731931580461039   0.8993565465052974   0.873612276320216   0.6641023513171929   0.8985866117995327   0.9488416160405383   0.8650812102986504   0.17440380184040785   0.33260524020991195   0.2536421899254926   0.05444919766029248   0.9727325085996703   0.60923822128941   0.5146356370203486   0.2402920414612218   0.9796891563655299   0.9197131523067379   0.8057692765453136   0.8679362499870272   0.03619933465056012   0.48232515401151227   0.23261011969704848   0.752413418769454   0.9981173304187507   0.9091319959654083   0.3332535731917511   0.878801142449238
0.33401497910155775   0.010545384165875629   0.3844119571512128   0.013719932150587678   0.15961117726114993   0.6779401439559637   0.1307697672257202   0.9592707344902952   0.18687866866147962   0.0687019226665538   0.6161341302053716   0.7189786930290734   0.20718951229594976   0.1489887703598159   0.810364853660058   0.8510424430420461   0.17099017764538965   0.6666636163483036   0.5777547339630095   0.09862902427259214   0.17287284722663895   0.7575316203828953   0.24450116077125836   0.21982788182335408   0.8388578681250812   0.7469862362170197   0.8600892036200456   0.20610794967276638   0.6792466908639313   0.06904609226105597   0.7293194363943254   0.2468372151824712   0.4923680222024517   0.00034416959450218106   0.11318530618895384   0.5278585221533978   0.2851785099065019   0.8513553992346863   0.30282045252889594   0.6768160791113517   0.11418833226111226   0.18469178288638266   0.7250657185658865   0.5781870548387595   0.9413154850344733   0.4271601625034874   0.48056455779462814   0.35835917301540543   0.1024576169093921   0.6801739262864677   0.6204753541745825   0.15225122334263905   0.42321092604546084   0.6111278340254117   0.8911559177802573   0.9054140081601678   0.9308429038430092   0.6107836644309095   0.7779706115913034   0.3775554860067701   0.6456643939365073   0.7594282651962232   0.47515015906240743   0.7007394068954184
0.5314760616753951   0.5747364823098405   0.7500844404965209   0.1225523520566589   0.5901605766409217   0.1475763198063532   0.2695198827018928   0.7641931790412535   0.4877029597315296   0.46740239351988555   0.6490445285273102   0.6119419556986144   0.06449203368606879   0.8562745594944738   0.7578886107470529   0.7065279475384466   0.1336491298430596   0.2454908950635643   0.9799179991557496   0.3289724615316765   0.48798473590655234   0.48606262986734106   0.5047678400933422   0.6282330546362581   0.9565086742311573   0.9113261475575005   0.7546833995968212   0.5056807025795992   0.36634809759023557   0.7637498277511473   0.4851635168949284   0.7414875235383457   0.8786451378587059   0.2963474342312618   0.8361189883676182   0.1295455678397313   0.8141531041726372   0.44007287473678797   0.07823037762056521   0.42301762030128476   0.6805039743295775   0.19458197967322366   0.09831237846481561   0.09404515876960826   0.19251923842302526   0.7085193498058826   0.5935445383714735   0.46581210413335017   0.23601056419186794   0.7971932022483821   0.8388611387746523   0.960131401553751   0.8696624666016324   0.03344337449723476   0.35369762187972387   0.21864387801540525   0.9910173287429265   0.737095940265973   0.5175786335121056   0.08909831017567393   0.17686422457028925   0.297023065529185   0.4393482558915404   0.6660806898743892
0.4963602502407117   0.10244108585596134   0.3410358774267248   0.5720355311047809   0.3038410118176864   0.39392173605007874   0.7474913390552513   0.10622342697143078   0.06783044762581847   0.5967285338016967   0.9086302002805992   0.1460920254176798   0.1981679810241861   0.5632851593044619   0.5549325784008753   0.9274481474022745   0.20715065228125967   0.826189219038489   0.037353944888769634   0.8383498372266006   0.03028642771097042   0.529166153509304   0.5980056889972292   0.17226914735221144   0.5339261774702587   0.4267250676533426   0.25696981157050436   0.6002336162474305   0.2300851656525723   0.03280333160326384   0.509478472515253   0.4940101892759997   0.16225471802675384   0.43607479780156716   0.6008482722346539   0.3479181638583199   0.9640867370025678   0.8727896384971052   0.04591569383377859   0.42047001645604537   0.756936084721308   0.046600419458616316   0.00856174894500895   0.5821201792294447   0.7266496570103377   0.5174342659493124   0.4105560599477798   0.4098510318772333   0.1927234795400789   0.0907091982959698   0.1535862483772754   0.8096174156298028   0.9626383138875066   0.057905866692705955   0.6441077758620224   0.3156072263538031   0.8003835958607528   0.6218310688911388   0.043259503627368516   0.9676890624954831   0.836296858858185   0.7490414303940335   0.9973438097935899   0.5472190460394378
0.07936077413687696   0.7024410109354172   0.988782060848581   0.965098866809993   0.3527111171265393   0.1850067449861048   0.5782260009008012   0.5552478349327598   0.1599876375864604   0.09429754669013503   0.42463975252352587   0.7456304193029569   0.1973493236989538   0.036391679997429066   0.7805319766615034   0.4300231929491538   0.39696572783820105   0.4145606111062903   0.7372724730341349   0.4623341304536706   0.560668868980016   0.6655191807122568   0.7399286632405451   0.9151150844142328   0.4813080948431391   0.9630781697768396   0.7511466023919641   0.9500162176042397   0.12859697771659975   0.7780714247907347   0.1729206014911628   0.39476838267148   0.9686093401301393   0.6837738781005996   0.7482808489676369   0.6491379633685231   0.7712600164311856   0.6473821981031707   0.9677488723061335   0.2191147704193693   0.37429428859298447   0.23282158699688035   0.23047639927199856   0.7567806399656987   0.8136254196129684   0.5673024062846236   0.4905477360314535   0.8416655555514658   0.3323173247698294   0.604224236507784   0.7394011336394894   0.8916493379472261   0.20372034705322964   0.8261528117170494   0.5664805321483267   0.49688095527574605   0.2351110069230903   0.14237893361644965   0.8181996831806897   0.8477429919072229   0.46385099049190476   0.49499673551327905   0.8504508108745562   0.6286282214878537
0.0895567018989203   0.2621751485163987   0.6199744116025576   0.8718475815221549   0.2759312822859519   0.6948727422317751   0.1294266755711041   0.030182025970689093   0.9436139575161224   0.09064850572399105   0.3900255419316146   0.138532688023463   0.7398936104628928   0.26449569400694173   0.8235450097832879   0.6416517327477169   0.5047826035398025   0.12211676039049203   0.00534532660259824   0.7939087408404939   0.040931613047897726   0.627120024877213   0.15489451572804203   0.1652805193526403   0.9513749111489774   0.3649448763608143   0.5349201041254844   0.29343293783048535   0.6754436288630256   0.6700721341290392   0.40549342855438025   0.26325091185979627   0.7318296713469031   0.5794236284050481   0.015467886622765653   0.12471822383633327   0.9919360608840103   0.3149279343981064   0.1919228768394777   0.4830664910886164   0.4871534573442078   0.19281117400761438   0.18657755023687947   0.6891577502481224   0.44622184429631007   0.5656911491304014   0.03168303450883743   0.5238772308954821   0.49484693314733263   0.20074627276958712   0.49676293038335306   0.23044429306499675   0.8194033042843071   0.5306741386405479   0.09126950182897277   0.9671933812052005   0.08757363293740396   0.9512505102354999   0.07580161520620711   0.8424751573688672   0.09563757205339367   0.6363225758373935   0.8838787383667294   0.35940866628025087
0.6084841147091858   0.4435114018297791   0.69730118812985   0.6702509160321285   0.1622622704128758   0.8778202526993777   0.6656181536210125   0.1463736851366464   0.6674153372655431   0.6770739799297906   0.16885522323765947   0.9159293920716496   0.8480120329812361   0.14639984128924263   0.0775857214086867   0.9487360108664491   0.7604384000438321   0.19514933105374277   0.0017841062024795868   0.10626085349758188   0.6648008279904385   0.5588267552163493   0.11790536783575017   0.746852187217331   0.05631671328125259   0.11531535338657023   0.42060417970590025   0.0766012711852025   0.8940544428683768   0.23749510068719254   0.7549860260848877   0.9302275860485562   0.22663910560283362   0.5604211207574019   0.5861308028472283   0.01429819397690651   0.37862707262159756   0.4140212794681593   0.5085450814385416   0.06556218311045739   0.6181886725777654   0.21887194841441657   0.506760975236062   0.9593013296128755   0.953387844587327   0.6600451931980672   0.3888556074003118   0.21244914239554452   0.8970711313060744   0.544729839811497   0.9682514276944115   0.135847871210342   0.003016688437697603   0.3072347391243045   0.2132654016095238   0.20562028516178588   0.776377582834864   0.7468136183669025   0.6271345987622956   0.19132209118487936   0.3977505102132664   0.3327923388987432   0.11858951732375399   0.12575990807442197
0.779561837635501   0.11392039048432662   0.611828542087692   0.16645857846154646   0.8261739930481741   0.45387519728625936   0.2229729346873802   0.954009436066002   0.9291028617420997   0.9091453574747623   0.25472150699296864   0.8181615648556599   0.926086173304402   0.6019106183504579   0.04145610538344482   0.6125412796938741   0.14970859046953805   0.8550969999835554   0.41432150662114925   0.42121918850899465   0.7519580802562716   0.5223046610848121   0.2957319892973953   0.2954592804345727   0.9723962426207706   0.40838427060048554   0.6839034472097033   0.12900070197302624   0.1462222495725966   0.9545090733142262   0.4609305125223231   0.1749912659070243   0.21711938783049697   0.04536371583946381   0.20620900552935445   0.35682970105136436   0.291033214526095   0.44345309748900597   0.16475290014590963   0.7442884213574903   0.1413246240565569   0.5883560975054506   0.7504313935247604   0.32306923284849565   0.3893665438002853   0.06605143642063846   0.4546994042273651   0.027609952413922962   0.4169703011795146   0.6576671658201529   0.7707959570176618   0.8986092504408967   0.270748051606918   0.7031580925059268   0.3098654444953387   0.7236179845338724   0.05362866377642103   0.657794376666463   0.1036564389659843   0.3667882834825081   0.7625954492503261   0.21434127917745702   0.9389035388200747   0.6224998621250177
0.6212708251937692   0.6259851816720065   0.1884721452953143   0.2994306292765221   0.2319042813934839   0.559933745251368   0.7337727410679492   0.27182067686259914   0.8149339802139692   0.902266579431215   0.9629767840502874   0.3732114264217024   0.5441859286070513   0.19910848692528824   0.6531113395549487   0.64959344188783   0.4905572648306302   0.5413141102588253   0.5494549005889644   0.2828051584053219   0.7279618155803042   0.32697283108136826   0.6105513617688897   0.6603052962803041   0.10669099038653497   0.7009876494093619   0.42207921647357544   0.36087466700378207   0.8747867089930511   0.1410539041579939   0.6883064754056262   0.08905399014118294   0.05985272877908182   0.2387873247267789   0.7253296913553388   0.7158425637194805   0.5156668001720306   0.03967883780149067   0.0722183518003901   0.06624912183165059   0.025109535341400365   0.4983647275426654   0.5227634512114258   0.7834439634263287   0.2971477197610962   0.17139189646129713   0.912212089442536   0.12313866714602455   0.19045672937456126   0.4704042470519353   0.4901328729689606   0.7622640001422425   0.31567002038151015   0.3293503428939414   0.8018263975633344   0.6732100100010595   0.25581729160242833   0.09056301816716246   0.07649670620799559   0.957367446281579   0.7401504914303978   0.0508841803656718   0.004278354407605494   0.8911183244499284
0.7150409560889974   0.5525194528230064   0.4815149031961798   0.10767436102359972   0.41789323632790115   0.38112755636170925   0.5693028137536438   0.9845356938775751   0.22743650695333992   0.910723309309774   0.07916994078468322   0.22227169373533268   0.9117664865718298   0.5813729664158326   0.27734354322134885   0.5490616837342731   0.6559491949694014   0.49080994824867014   0.20084683701335324   0.5916942374526941   0.9157987035390036   0.43992576788299836   0.19656848260574775   0.7005759130027657   0.20075774745000624   0.8874063150599919   0.7150535794095679   0.592901551979166   0.7828645111221051   0.5062787586982826   0.14575076565592418   0.6083658581015908   0.5554280041687651   0.5955554493885087   0.06658082487124095   0.38609416436625815   0.6436615175969354   0.014182482972676089   0.7892372816498922   0.837032480631985   0.987712322627534   0.5233725347240059   0.5883904446365389   0.2453382431792909   0.07191361908853033   0.08344676684100759   0.3918219620307911   0.5447623301765252   0.871155871638524   0.19604045178101562   0.6767683826212232   0.9518607781973591   0.088291360516419   0.6897616930827329   0.531017616965299   0.3434949200957683   0.5328633563476538   0.09420624369422423   0.4644367920940581   0.9574007557295101   0.8892018387507185   0.08002376072154814   0.6751995104441659   0.12036827509752511
0.9014895161231845   0.5566512259975422   0.08680906580762705   0.8750300319182343   0.8295758970346542   0.47320445915653464   0.6949871037768359   0.33026770174170905   0.9584200253961301   0.277164007375519   0.018218721155612724   0.37840692354434985   0.8701286648797111   0.5874023142927861   0.4872011041903137   0.034912003448581544   0.3372653085320572   0.4931960705985618   0.022764312096255658   0.07751124771907139   0.44806346978133876   0.4131723098770137   0.34756480165208975   0.9571429726215462   0.5465739536581543   0.8565210838794715   0.26075573584446265   0.08211294070331207   0.7169980566235001   0.3833166247229368   0.5657686320676267   0.751845238961603   0.75857803122737   0.10615261734741785   0.547549910912014   0.3734383154172532   0.8884493663476589   0.5187503030546318   0.060348806721700336   0.33852631196867167   0.5511840578156016   0.02555423245606997   0.03758449462544468   0.26101506424960025   0.10312058803426294   0.6123819225790563   0.690019692973355   0.30387209162805395   0.5565466343761087   0.7558608386995849   0.42926395712889226   0.22175915092474188   0.8395485777526086   0.372544213976648   0.8634953250612655   0.46991391196313886   0.08097054652523861   0.2663915966292302   0.3159454141492515   0.09647559654588565   0.1925211801775797   0.7476412935745984   0.25559660742755114   0.757949284577214
0.641337122361978   0.7220870611185284   0.21801211280210644   0.49693422032761375   0.538216534327715   0.1097051385394721   0.5279924198287514   0.19306212869955977   0.9816698999516064   0.35384429983988724   0.09872846269985922   0.9713029777748179   0.14212132219899776   0.9813000858632392   0.23523313763859371   0.5013890658116791   0.06115077567375915   0.7149084892340091   0.9192877234893423   0.4049134692657934   0.8686295954961795   0.9672671956594108   0.6636911160617911   0.6469641846885794   0.22729247313420148   0.24518013454088236   0.4456790032596847   0.15002996436096563   0.6890759388064864   0.13547499600141027   0.9176865834309332   0.9569678356614059   0.7074060388548801   0.781630696161523   0.818958120731074   0.985664857886588   0.5652847166558823   0.8003306102982837   0.5837249830924802   0.48427579207490895   0.5041339409821232   0.0854221210642746   0.664437259603138   0.07936232280911555   0.6355043454859437   0.11815492540486384   0.0007461435413468715   0.4323981381205362   0.4082118723517422   0.8729747908639814   0.5550671402816622   0.2823681737595705   0.7191359335452558   0.7374997948625712   0.637380556850729   0.32540033809816465   0.011729894690375707   0.9558690987010482   0.818422436119655   0.3397354802115767   0.44644517803449335   0.1555384884027645   0.23469745302717474   0.8554596881366677
0.9423112370523702   0.07011636733848989   0.5702601934240367   0.7760973653275522   0.3068068915664265   0.9519614419336261   0.5695140498826898   0.34369922720701607   0.8985950192146842   0.07898665106964456   0.014446909601027664   0.06133105344744553   0.17945908566942845   0.34148685620707336   0.3770663527502987   0.7359307153492809   0.16772919097905276   0.3856177575060251   0.5586439166306437   0.39619523513770416   0.7212840129445593   0.23007926910326063   0.32394646360346896   0.5407355470010364   0.7789727758921892   0.15996290176477074   0.7536862701794322   0.7646381816734842   0.4721658843257627   0.20800145983114468   0.1841722202967424   0.4209389544664681   0.5735708651110785   0.12901480876150012   0.16972531069571475   0.35960790101902257   0.39411177944165   0.7875279525544268   0.7926589579454161   0.6236771856697417   0.22638258846259723   0.4019101950484017   0.23401504131477235   0.22748195053203757   0.5050985755180378   0.17183092594514107   0.9100685777113033   0.6867464035310011   0.7261257996258487   0.011868024180370331   0.15638230753187113   0.922108221857517   0.253959915300086   0.8038665643492257   0.9722100872351287   0.5011692673910488   0.6803890501890075   0.6748517555877255   0.802484776539414   0.1415613663720263   0.28627727074735754   0.8873238030332987   0.009825818593997906   0.5178841807022846
0.0598946822847603   0.485413607984897   0.7758107772792255   0.29040223017024697   0.5547961067667224   0.313582682039756   0.8657421995679222   0.6036558266392458   0.8286703071408738   0.3017146578593856   0.709359892036051   0.6815476047817288   0.5747103918407878   0.49784809351016   0.7371498048009223   0.18037833739067993   0.8943213416517802   0.8229963379224345   0.9346650282615083   0.03881697101865364   0.6080440709044227   0.9356725348891358   0.9248392096675104   0.5209327903163691   0.5481493886196624   0.45025892690423874   0.14902843238828486   0.2305305601461221   0.99335328185294   0.1366762448644828   0.28328623282036275   0.6268747335068763   0.16468297471206622   0.8349615870050972   0.5739263407843117   0.9453271287251476   0.5899725828712784   0.33711349349493713   0.8367765359833894   0.7649487913344676   0.6956512412194982   0.5141171555725027   0.9021115077218811   0.7261318203158139   0.08760717031507545   0.5784446206833669   0.9772722980543707   0.20519902999944487   0.539457781695413   0.12818569377912814   0.8282438656660858   0.9746684698533228   0.5461044998424731   0.9915094489146453   0.5449576328457231   0.34779373634644645   0.38142152513040684   0.15654786190954822   0.9710312920614114   0.40246660762129893   0.7914489422591284   0.819434368414611   0.13425475607802193   0.6375178162868314
0.09579770103963026   0.3053172128421084   0.23214324835614084   0.9113859959710173   0.008190530724554803   0.7268725921587414   0.25487095030177015   0.7061869659715725   0.46873274902914175   0.5986868983796133   0.42662708463568433   0.7315184961182497   0.9226282491866687   0.607177449464968   0.8816694517899613   0.3837247597718033   0.5412067240562618   0.45062958755541976   0.9106381597285499   0.9812581521505044   0.7497577817971334   0.6311952191408087   0.7763834036505279   0.3437403358636731   0.6539600807575031   0.3258780062987003   0.5442401552943871   0.4323543398926557   0.6457695500329483   0.5990054141399588   0.289369204992617   0.7261673739210832   0.1770368010038066   0.00031851576034545555   0.8627421203569327   0.9946488778028335   0.2544085518171379   0.3931410662953775   0.9810726685669714   0.6109241180310302   0.713201827760876   0.9425114787399577   0.07043450883842149   0.6296659658805258   0.9634440459637427   0.311316259599149   0.2940511051878935   0.2859256300168528   0.30948396520623944   0.9854382533004487   0.7498109498935064   0.8535712901241971   0.6637144151732911   0.38643283916048987   0.46044174490088946   0.1274039162031138   0.4866776141694845   0.3861143234001444   0.5976996245439568   0.1327550384002803   0.2322690623523466   0.9929732571047669   0.6166269559769854   0.52183092036925
0.5190672345914705   0.05046177836480925   0.546192447138564   0.8921649544887242   0.555623188627728   0.7391455187656603   0.2521413419506704   0.6062393244718715   0.24613922342148847   0.7537072654652116   0.502330392057164   0.7526680343476745   0.5824248082481974   0.3672744263047217   0.04188864715627452   0.6252641181445606   0.09574719407871289   0.9811601029045773   0.44418902261231774   0.4925090797442803   0.8634781317263663   0.9881868457998103   0.8275620666353323   0.9706781593750302   0.34441089713489575   0.9377250674350011   0.2813696194967684   0.07851320488630595   0.7887877085071678   0.19857954866934083   0.029228277546098035   0.47227388041443447   0.5426484850856793   0.44487228320412925   0.5268978854889341   0.71960584606676   0.960223676837482   0.07759785689940754   0.4850092383326596   0.0943417279221994   0.8644764827587691   0.09643775399483026   0.04082021572034183   0.6018326481779191   0.0009983510324027766   0.10825090819501992   0.2132581490850095   0.6311544888028889   0.6565874538975071   0.17052584076001884   0.9318885295882411   0.552641283916583   0.8677997453903392   0.971946292090678   0.9026602520421431   0.08036740350214851   0.32515126030465985   0.5270740088865488   0.375762366553209   0.3607615574353885   0.3649275834671779   0.4494761519871412   0.8907531282205494   0.2664198295131891
0.5004511007084088   0.35303839799231096   0.8499329125002076   0.66458718133527   0.49945274967600606   0.24478748979729104   0.6366747634151981   0.03343269253238108   0.842865295778499   0.0742616490372722   0.704786233826957   0.4807914086157981   0.9750655503881598   0.10231535694659419   0.802125981784814   0.4004240051136496   0.6499142900835   0.5752413480600455   0.42636361523160493   0.03966244767826111   0.284986706616322   0.1257651960729042   0.5356104870110555   0.773242618165072   0.7845356059079132   0.7727267980805933   0.6856775745108479   0.10865543682980204   0.2850828562319071   0.5279393082833023   0.0490028110956498   0.07522274429742097   0.4422175604534081   0.45367765924603004   0.3442165772686928   0.5944313356816229   0.46715201006524826   0.3513623022994358   0.5420905954838788   0.19400733056797326   0.8172377199817483   0.7761209542393904   0.11572698025227396   0.15434488288971215   0.5322510133654264   0.6503557581664862   0.5801164932412185   0.3811022647246401   0.7477154074575131   0.8776289600858929   0.8944389187303705   0.2724468278948381   0.462632551225606   0.3496896518025907   0.8454361076347208   0.1972240835974171   0.020414990772197914   0.8960119925565606   0.501219530366028   0.6027927479157943   0.5532629807069497   0.5446496902571248   0.959128934882149   0.408785417347821
0.7360252607252014   0.7685287360177344   0.8434019546298751   0.2544405344581088   0.20377424735977503   0.11817297785124826   0.26328546138865666   0.8733382697334687   0.4560588399022619   0.24054401776535533   0.3688465426582861   0.6008914418386306   0.9934262886766559   0.8908543659627647   0.5234104350235653   0.4036673582412136   0.973011297904458   0.994842373406204   0.022190904657537397   0.8008746103254193   0.4197483171975084   0.4501926831490792   0.06306196977538835   0.3920891929775983   0.683723056472307   0.6816639471313447   0.21966001514551325   0.1376486585194895   0.479948809112532   0.5634909692800965   0.9563745537568565   0.26431038878602076   0.02388996921027009   0.3229469515147411   0.5875280110985704   0.6634189469473901   0.030463680533614174   0.43209258555197644   0.06411757607500516   0.25975158870617654   0.05745238262915617   0.4372502121457725   0.04192667141746776   0.45887697838075725   0.6377040654316478   0.9870575289966933   0.9788647016420794   0.0667877854031589   0.9539810089593408   0.3053935818653486   0.7592046864965661   0.9291391268836694   0.4740321998468088   0.7419026125852521   0.8028301327397096   0.6648287380976486   0.4501422306365387   0.41895566107051097   0.21530212164113907   0.001409791150258549   0.41967855010292454   0.9868630755185345   0.15118454556613392   0.741658202444082
0.36222616747376835   0.549612863372762   0.10925787414866617   0.2827812240633248   0.7245221020421205   0.5625553343760687   0.13039317250658675   0.21599343866016588   0.7705410930827797   0.2571617525107202   0.3711884860100206   0.28685431177649645   0.29650889323597096   0.5152591399254681   0.568358353270311   0.6220255736788478   0.8463666625994323   0.0963034788549571   0.35305623162917193   0.6206157825285893   0.4266881124965078   0.10944040333642259   0.201871686063038   0.8789575800845072   0.06446194502273943   0.5598275399636605   0.09261381191437182   0.5961763560211825   0.3399398429806189   0.9972722055875918   0.962220639407785   0.3801829173610166   0.5693987498978391   0.7401104530768716   0.5910321533977645   0.09332860558452016   0.27288985666186816   0.22485131315140353   0.022673800127453493   0.47130303190567235   0.4265231940624359   0.12854783429644642   0.6696175684982816   0.8506872493770832   0.9998350815659282   0.019107430960023822   0.4677458824352436   0.9717296692925759   0.9353731365431887   0.4592798909963633   0.3751320705208718   0.3755533132713934   0.5954332935625698   0.4620076854087715   0.41291143111308676   0.9953703959103768   0.026034543664730663   0.7218972323318998   0.8218792777153222   0.9020417903258566   0.7531446870028625   0.49704591918049634   0.7992054775878688   0.4307387584201843
0.3266214929404266   0.36849808488404995   0.12958790908958717   0.5800515090431011   0.3267864113744985   0.34939065392402613   0.6618420266543436   0.6083218397505252   0.3914132748313098   0.8901107629276629   0.2867099561334718   0.23276852647913182   0.7959799812687399   0.4281030775188914   0.873798525020385   0.23739813056875503   0.7699454376040092   0.7062058451869915   0.051919247305062796   0.3353563402428984   0.016800750601146792   0.2091599260064951   0.25271376971719406   0.9046175818227141   0.6901792576607202   0.8406618411224451   0.12312586062760687   0.324566072779613   0.36339284628622176   0.491271187198419   0.46128383397326334   0.7162442330290878   0.971979571454912   0.6011604242707562   0.17457387783979153   0.483475706549956   0.17599959018617203   0.17305734675186482   0.3007753528194065   0.24607757598120092   0.40605415258216276   0.4668515015648734   0.2488561055143437   0.9107212357383025   0.389253401981016   0.2576915755583783   0.9961423357971496   0.006103653915588378   0.6990741443202958   0.4170297344359331   0.8730164751695427   0.6815375811359754   0.33568129803407404   0.925758547237514   0.41173264119627945   0.9652933481068876   0.36370172657916205   0.32459812296675794   0.23715876335648794   0.48181764155693163   0.18770213639299   0.1515407762148931   0.9363834105370814   0.23574006557573068
0.7816479838108272   0.6846892746500197   0.6875273050227377   0.3250188298374282   0.3923945818298113   0.4269976990916414   0.6913849692255881   0.3189151759218398   0.6933204375095156   0.009967964655708322   0.8183684940560453   0.6373775947858644   0.35763913947544146   0.08420941741819422   0.40663585285976583   0.6720842466789768   0.9939374128962795   0.7596112944514363   0.1694770895032779   0.19026660512204524   0.8062352765032894   0.6080705182365432   0.23309367896619645   0.9545265395463145   0.02458729269246221   0.9233812435865235   0.5455663739434587   0.6295077097088864   0.6321927108626509   0.49638354449488203   0.8541814047178706   0.31059253378704654   0.9388722733531354   0.4864155798391737   0.035812910661825355   0.6732149390011821   0.5812331338776939   0.4022061624209795   0.6291770578020596   0.001130692322205273   0.5872957209814145   0.6425948679695432   0.4596999682987816   0.81086408720016   0.7810604444781251   0.03452434973299999   0.22660628933258517   0.8563375476538455   0.7564731517856629   0.11114310614647652   0.6810399153891264   0.22682983794495915   0.12428044092301192   0.6147595616515945   0.8268585106712558   0.9162373041579126   0.1854081675698765   0.12834398181242077   0.7910456000094305   0.24302236515673042   0.6041750336921825   0.7261378193914413   0.16186854220737093   0.24189167283452515
0.01687931271076801   0.08354295142189808   0.7021685739085893   0.4310275856343651   0.23581886823264295   0.049018601688898086   0.4755622845760041   0.5746900379805197   0.4793457164469801   0.9378754955424216   0.7945223691868777   0.3478602000355605   0.35506527552396816   0.3231159338908271   0.9676638585156219   0.4316228958776479   0.16965710795409167   0.19477195207840634   0.1766182585061914   0.1886005307209175   0.5654820742619091   0.468634132686965   0.014749716298820466   0.9467088578863924   0.5486027615511411   0.385091181265067   0.31258114239023116   0.5156812722520272   0.31278389331849815   0.3360725795761689   0.837018857814227   0.9409912342715075   0.8334381768715181   0.3981970840337473   0.04249648862734942   0.5931310342359472   0.47837290134754995   0.0750811501429202   0.07483263011172758   0.16150813835829916   0.3087157933934583   0.8803091980645139   0.8982143716055362   0.9729076076373817   0.7432337191315491   0.41167506537754883   0.8834646553067157   0.026198749750989334   0.19463095758040805   0.026583884112481863   0.5708835129164845   0.5105174774989621   0.8818470642619098   0.690511304536313   0.7338646551022575   0.5695262432274545   0.048408887390391765   0.29231422050256567   0.6913681664749081   0.9763952089915074   0.5700359860428418   0.21723307035964548   0.6165355363631805   0.8148870706332082
0.2613201926493835   0.3369238722951316   0.7183211647576443   0.8419794629958266   0.5180864735178343   0.9252488069175828   0.8348565094509286   0.8157807132448373   0.3234555159374263   0.8986649228051009   0.263972996534444   0.3052632357458751   0.44160845167551643   0.20815361826878792   0.5301083414321865   0.7357369925184206   0.39319956428512465   0.9158393977662223   0.8387401749572785   0.7593417835269132   0.8231635782422828   0.6986063274065768   0.22220463859409803   0.944454712893705   0.5618433855928994   0.36168245511144514   0.5038834738364537   0.10247524989787836   0.04375691207506499   0.4364336481938624   0.6690269643855252   0.2866945366530411   0.7203013961376387   0.5377687253887614   0.40505396785108116   0.981431300907166   0.2786929444621223   0.3296151071199735   0.8749456264188946   0.2456943083887454   0.8854933801769976   0.41377570935375124   0.03620545146161614   0.4863525248618322   0.06232980193471479   0.7151693819471745   0.8140008128675181   0.5418978119681273   0.5004864163418155   0.35348692683572935   0.31011733903106437   0.43942256207024893   0.45672950426675046   0.917053278641867   0.6410903746455392   0.1527280254172078   0.7364281081291117   0.37928455325310556   0.23603640679445795   0.17129672451004183   0.45773516366698946   0.049669446133132046   0.3610907803755633   0.9256024161212965
0.5722417834899919   0.6358937367793808   0.32488532891394717   0.4392498912594642   0.5099119815552771   0.9207243548322063   0.510884516046429   0.8973520792913369   0.009425565213461587   0.5672374279964769   0.20076717701536473   0.45792951722108793   0.5526960609467111   0.6501841493546099   0.5596768023698255   0.3052014918038801   0.8162679528175993   0.2708995961015044   0.3236403955753676   0.1339047672938383   0.3585327891506099   0.22123014996837234   0.9625496151998043   0.2083023511725419   0.786291005660618   0.5853364131889915   0.6376642862858571   0.7690524599130777   0.27637902410534104   0.6646120583567853   0.12677977023942805   0.8717003806217408   0.26695345889187944   0.09737463036030834   0.9260125932240634   0.4137708634006529   0.7142573979451683   0.4471904810056984   0.36633579085423773   0.10856937159677274   0.897989445127569   0.17629088490419403   0.042695395278870125   0.9746646043029344   0.539456655976959   0.9550607349358217   0.08014578007906584   0.7663622531303925   0.753165650316341   0.3697243217468302   0.4424814937932087   0.9973097932173148   0.47678662621099993   0.7051122633900448   0.3157017235537807   0.12560941259557407   0.20983316731912052   0.6077376330297365   0.38968913032971736   0.7118385491949212   0.4955757693739522   0.16054715202403813   0.02335333947547961   0.6032691775981485
0.5975863242463832   0.9842562671198442   0.9806579441966095   0.628604573295214   0.058129668269424235   0.02919553218402241   0.9005121641175436   0.8622423201648215   0.30496401795308326   0.6594712104371923   0.4580306703243349   0.8649325269475066   0.8281773917420833   0.9543589470471474   0.14232894677055427   0.7393231143519325   0.6183442244229628   0.3466213140174108   0.7526398164408369   0.027484565157011316   0.12276845504901057   0.1860741619933727   0.7292864769653573   0.42421538755886284   0.5251821308026273   0.20181789487352858   0.7486285327687479   0.7956108142636489   0.46705246253320304   0.17262236268950618   0.8481163686512042   0.9333684940988274   0.16208844458011978   0.5131511522523139   0.39008569832686923   0.06843596715132083   0.33391105283803646   0.5587922052051665   0.24775675155631496   0.32911285279938834   0.7155668284150737   0.2121708911877557   0.49511693511547805   0.301628287642377   0.5927983733660631   0.026096729194383005   0.7658304581501207   0.8774129000835141   0.06761624256343585   0.8242788343208545   0.01720192538137294   0.08180208581986528   0.6005637800302328   0.6516564716313482   0.16908555673016878   0.14843359172103787   0.438475335450113   0.13850531937903435   0.7789998584032995   0.07999762456971704   0.10456428261207652   0.5797131141738678   0.5312431068469846   0.7508847717703288
0.3889974541970028   0.3675422229861121   0.03612617173150654   0.4492564841279517   0.7961990808309397   0.3414454937917291   0.27029571358138577   0.5718435840444376   0.7285828382675038   0.5171666594708747   0.2530937882000128   0.49004149822457227   0.12801905823727106   0.8655101878395264   0.08400823146984407   0.3416079065035344   0.689543722787158   0.7270048684604921   0.3050083730665445   0.26161028193381736   0.5849794401750815   0.14729175428662428   0.7737652662195599   0.5107255101634887   0.19598198597807873   0.7797495313005122   0.7376390944880534   0.06146902603553695   0.39978290514713904   0.43830403750878305   0.4673433809066676   0.48962544199109936   0.6712000668796352   0.9211373780379084   0.21424959270665472   0.999583943766527   0.5431810086423642   0.055627190198381964   0.13024136123681065   0.6579760372629927   0.853637285855206   0.32862232173788986   0.8252329881702661   0.3963657553291753   0.2686578456801246   0.1813305674512656   0.051467721950706244   0.8856402451656866   0.07267585970204585   0.4015810361507534   0.3138286274626529   0.8241712191301497   0.6728929545549068   0.9632769986419704   0.8464852465559853   0.3345457771390503   0.0016928876752716144   0.042139620604061956   0.6322356538493306   0.3349618333725232   0.45851187903290747   0.98651243040568   0.5019942926125199   0.6769857961095306
0.6048745931777014   0.6578901086677901   0.6767613044422537   0.28062004078035524   0.3362167474975768   0.4765595412165245   0.6252935824915475   0.3949797956146686   0.263540887795531   0.0749785050657711   0.3114649550288946   0.570808576484519   0.5906479332406241   0.11170150642380075   0.4649797084729093   0.23626279934546862   0.5889550455653525   0.0695618858197388   0.8327440546235788   0.9013009659729454   0.1304431665324451   0.0830494554140588   0.3307497620110589   0.22431516986341488   0.5255685733547437   0.4251593467462687   0.6539884575688052   0.9436951290830596   0.1893518258571669   0.9485998055297442   0.02869487507725767   0.548715333468391   0.925810938061636   0.873621300463973   0.7172299200483631   0.9779067569838721   0.33516300482101175   0.7619197940401723   0.25225021157545374   0.7416439576384034   0.7462079592556592   0.6923579082204335   0.41950615695187493   0.840342991665458   0.6157647927232142   0.6093084528063747   0.08875639494081607   0.6160278218020432   0.0901962193684704   0.18414910606010604   0.4347679373720109   0.6723326927189835   0.9008443935113035   0.23554930053036188   0.40607306229475326   0.12361735925059253   0.9750334554496676   0.3619280000663888   0.6888431422463902   0.14571060226672047   0.6398704506286559   0.6000082060262165   0.43659293067093646   0.40406664462831704
0.8936624913729967   0.907650297805783   0.017086773719061508   0.563723652962859   0.27789769864978253   0.2983418449994083   0.9283303787782454   0.9476958311608159   0.18770147928131214   0.11419273893930224   0.4935624414062345   0.27536313844183236   0.2868570857700086   0.8786434384089403   0.08748937911148129   0.15174577919123983   0.31182363032034105   0.5167154383425515   0.3986462368650911   0.006035176924519344   0.6719531796916851   0.916707232316335   0.9620533061941546   0.6019685322962023   0.7782906883186885   0.009056934510552006   0.9449665324750931   0.038244879333343265   0.5003929896689059   0.7107150895111437   0.0166361536968477   0.09054904817252739   0.3126915103875938   0.5965223505718416   0.5230737122906132   0.815185909730695   0.025834424617585148   0.7178789121629011   0.43558433317913187   0.6634401305394552   0.7140107942972441   0.20116347382034963   0.036938096314040755   0.6574049536149359   0.042057614605558964   0.2844562415040146   0.07488479011988611   0.055436421318733574   0.2637669262868705   0.2753993069934626   0.12991825764479298   0.017191541985390305   0.7633739366179646   0.5646842174823189   0.11328210394794527   0.9266424938128629   0.45068242623037075   0.9681618669104773   0.5902083916573321   0.1114565840821679   0.42484800161278563   0.2502829547475762   0.15462405847820024   0.4480164535427127
0.7108372073155415   0.04911948092722661   0.11768596216415948   0.7906114999277768   0.6687795927099826   0.764663239423212   0.042801172044273375   0.7351750786090432   0.40501266642311207   0.48926393242974936   0.9128829143994804   0.7179835366236529   0.6416387298051475   0.9245797149474305   0.7996008104515351   0.79134104281079   0.19095630357477675   0.9564178480369531   0.20939241879420303   0.6798844587286221   0.7661083019619911   0.7061348932893768   0.05476836031600278   0.23186800518590944   0.05527109464644962   0.6570154123621502   0.9370823981518432   0.44125650525813265   0.3864915019364671   0.8923521729389383   0.8942812261075699   0.7060814266490893   0.981478835513355   0.4030882405091889   0.9813983117080896   0.9880978900254365   0.3398401057082075   0.47850852556175844   0.1817975012565544   0.19675684721464648   0.14888380213343078   0.5220906775248053   0.9724050824623514   0.5168723884860243   0.38277550017143963   0.8159557842354285   0.9176367221463486   0.2850043833001149   0.32750440552499005   0.15894037187327822   0.9805543239945053   0.8437478780419823   0.941012903588523   0.26658819893433994   0.08627309788693537   0.13766645139289288   0.959534068075168   0.863499958425151   0.10487478617884584   0.14956856136745642   0.6196939623669604   0.38499143286339266   0.9230772849222915   0.95281171415281
0.4708101602335296   0.8629007553385873   0.9506722024599401   0.43593932566678556   0.08803466006208996   0.046944971103158845   0.03303548031359149   0.15093494236667068   0.7605302545370999   0.8880045992298806   0.0524811563190862   0.3071870643246884   0.819517350948577   0.6214164002955407   0.9662080584321509   0.16952061293179552   0.8599832828734091   0.7579164418703896   0.861333272253305   0.01995205156433912   0.2402893205064487   0.372925009006997   0.9382559873310136   0.06714033741152918   0.7694791602729191   0.5100242536684096   0.9875837848710735   0.6312010117447436   0.6814445002108291   0.4630792825652508   0.954548304557482   0.4802660693780729   0.9209142456737291   0.5750746833353703   0.9020671482383957   0.17307900505338453   0.1013968947251522   0.9536582830398296   0.9358590898062449   0.003558392121589011   0.24141361185174315   0.1957418411694399   0.07452581755293994   0.9836063405572499   0.0011242913452944603   0.822816832162443   0.1362698302219264   0.9164660031457207   0.2316451310723754   0.31279257849403325   0.14868604535085295   0.2852649914009771   0.5502006308615462   0.8497132959287824   0.19413774079337098   0.8049989220229041   0.6292863851878171   0.2746386125934122   0.2920705925549752   0.6319199169695197   0.5278894904626649   0.3209803295535827   0.35621150274873026   0.6283615248479306
0.2864758786109218   0.12523848838414275   0.28168568519579035   0.6447551842906807   0.2853515872656273   0.3024216562216998   0.14541585497386394   0.72828918114496   0.0537064561932519   0.9896290777276666   0.996729809623011   0.44302418974398294   0.5035058253317056   0.13991578179888414   0.8025920688296401   0.6380252677210787   0.8742194401438885   0.8652771692054719   0.5105214762746648   0.006105350751559118   0.3463299496812236   0.5442968396518892   0.15430997352593456   0.3777438259036285   0.05985407107030186   0.41905835126774654   0.8726242883301443   0.7329886416129477   0.7745024838046746   0.11663669504604669   0.7272084333562803   0.004699460467987718   0.7207960276114227   0.12700761731838012   0.7304786237332692   0.5616752707240048   0.21729020227971707   0.987091835519496   0.9278865549036293   0.923650003002926   0.34307076213582854   0.12181466631402402   0.4173650786289644   0.9175446522513669   0.9967408124546049   0.5775178266621347   0.2630551051030298   0.5398008263477384   0.9368867413843031   0.15845947539438823   0.3904308167728856   0.8068121847347907   0.1623842575796285   0.04182278034834152   0.6632223834166053   0.8021127242668029   0.4415882299682058   0.9148151630299614   0.9327437596833361   0.24043745354279816   0.22429802768848875   0.9277233275104654   0.004857204779706855   0.3167874505398721
0.8812272655526602   0.8059086611964414   0.5874921261507424   0.39924279828850523   0.8844864530980553   0.22839083453430667   0.32443702104771266   0.8594419719407668   0.9475997117137522   0.06993135913991844   0.9340062042748271   0.052629787205976136   0.7852154541341237   0.028108578791576917   0.27078382085822167   0.2505170629391732   0.3436272241659179   0.11329341576161553   0.3380400611748856   0.010079609396375018   0.11932919647742916   0.1855700882511501   0.33318285639517875   0.6932921588565029   0.23810193092476895   0.3796614270547087   0.7456907302444362   0.29404936056799763   0.35361547782671365   0.15127059252040204   0.4212537091967236   0.43460738862723086   0.4060157661129615   0.0813392333804836   0.4872475049218966   0.3819776014212547   0.6208003119788377   0.05323065458890669   0.21646368406367494   0.13146053848208153   0.27717308781291977   0.9399372388272912   0.8784236228887894   0.12138092908570652   0.15784389133549065   0.754367150576141   0.5452407664936106   0.42808877022920366   0.9197419604107216   0.3747057235214324   0.7995500362491743   0.13403940966120598   0.566126482584008   0.22343513100103032   0.3782963270524507   0.6994320210339752   0.16011071647104658   0.14209589762054672   0.891048822130554   0.3174544196127204   0.5393104044922089   0.08886524303164003   0.6745851380668791   0.18599388113063886
0.2621373166792891   0.14892800420434887   0.7961615151780898   0.06461295204493235   0.10429342534379843   0.3945608536282078   0.25092074868447917   0.6365241818157287   0.18455146493307675   0.01985513010677544   0.4513707124353048   0.5024847721545227   0.6184249823490687   0.7964199991057451   0.0730743853828541   0.8030527511205476   0.45831426587802215   0.6543241014851984   0.18202556325230002   0.48559833150782716   0.9190038613858132   0.5654588584535584   0.5074404251854209   0.2996044503771883   0.6568665447065243   0.4165308542492095   0.7112789100073311   0.23499149833225597   0.5525731193627258   0.02197000062100168   0.46035816132285196   0.5984673165165273   0.36802165442964907   0.0021148705142262393   0.008987448887547147   0.09598254436200453   0.7495966720805803   0.2056948714084811   0.935913063504693   0.2929297932414569   0.2912824062025582   0.5513707699232827   0.753887500252393   0.8073314617336297   0.3722785448167449   0.9859119114697243   0.2464470750669721   0.5077270113564414   0.7154120001102207   0.5693810572205149   0.535168165059641   0.27273551302418547   0.16283888074749484   0.5474110565995132   0.07481000373678905   0.6742681965076582   0.7948172263178458   0.545296186085287   0.0658225548492419   0.5782856521456536   0.045220554237265405   0.3396013146768058   0.12990949134454885   0.28535585890419674
0.7539381480347072   0.788230544753523   0.37602199109215584   0.478024397170567   0.38165960321796233   0.8023186332837987   0.12957491602518373   0.9702973858141256   0.6662476031077417   0.23293757606328386   0.5944067509655427   0.6975618727899402   0.5034087223602468   0.6855265194637706   0.5195967472287537   0.02329367628228197   0.708591496042401   0.1402303333784837   0.4537741923795118   0.4450080241366283   0.6633709418051357   0.8006290187016779   0.3238647010349629   0.15965216523243156   0.9094327937704284   0.012398473948154758   0.9478427099428071   0.6816277680618645   0.5277731905524661   0.210079840664356   0.8182677939176234   0.7113303822477389   0.8615255874447245   0.9771422646010721   0.22386104295208065   0.013768509457798757   0.35811686508447765   0.2916157451373015   0.7042642957233269   0.9904748331755168   0.6495253690420766   0.15138541175881778   0.2504901033438152   0.5454668090388884   0.9861544272369409   0.3507563930571399   0.9266254023088523   0.3858146438064569   0.07672163346651248   0.33835791910898516   0.9787826923660452   0.7041868757445924   0.5489484429140463   0.12827807844462916   0.16051489844842187   0.9928564934968535   0.6874228554693219   0.15113581384355698   0.9366538554963413   0.9790879840390547   0.32930599038484426   0.8595200687062555   0.23238955977301426   0.988613150863538
0.6797806213427676   0.7081346569474377   0.9818994564291991   0.44314634182464946   0.6936261941058267   0.3573782638902978   0.05527405412034677   0.05733169801819252   0.6169045606393142   0.019020344781312617   0.07649136175430155   0.3531448222736001   0.0679561177252679   0.8907422663366835   0.9159764633058797   0.3602883287767466   0.380533262255946   0.7396064524931265   0.9793226078095385   0.3812003447376919   0.05122727187110177   0.880086383786871   0.7469330480365242   0.3925871938741539   0.3714466505283341   0.17195172683943327   0.7650335916073251   0.9494408520495045   0.6778204564225073   0.8145734629491355   0.7097595374869784   0.892109154031312   0.060915895783193126   0.7955531181678228   0.6332681757326768   0.5389643317577119   0.9929597780579252   0.9048108518311394   0.7172917124267971   0.17867600298096525   0.6124265158019793   0.16520439933801292   0.7379691046172587   0.7974756582432734   0.5611992439308774   0.28511801555114197   0.9910360565807345   0.4048884643691194   0.18975259340254333   0.11316628871170868   0.22600246497340937   0.45544761231961495   0.5119321369800359   0.2985928257625732   0.516242927486431   0.563338458288303   0.4510162411968428   0.5030397075947504   0.8829747517537542   0.024374126530591095   0.4580564631389176   0.598228855763611   0.16568303932695702   0.8456981235496258
0.8456299473369384   0.433024456425598   0.4277139347096984   0.0482224653063525   0.28443070340606097   0.14790644087445606   0.43667787812896386   0.6433340009372331   0.09467811000351761   0.03474015216274738   0.2106754131555545   0.18788638861761817   0.5827459730234816   0.7361473264001742   0.6944324856691235   0.6245479303293152   0.13172973182663883   0.23310761880542386   0.8114577339153694   0.6001738037987241   0.6736732686877213   0.6348787630418129   0.6457746945884123   0.7544756802490983   0.8280433213507828   0.20185430661621495   0.21806075987871396   0.7062532149427457   0.5436126179447219   0.05394786574175888   0.7813828817497501   0.06291921400551267   0.44893450794120426   0.019207713579011496   0.5707074685941956   0.8750328253878945   0.8661885349177226   0.2830603871788373   0.8762749829250721   0.2504848950585793   0.7344588030910838   0.049952768373413434   0.06481724900970276   0.6503110912598552   0.060785534403362554   0.4150740053316005   0.41904255442129046   0.8958354110107569   0.23274221305257972   0.21321969871538557   0.2009817945425765   0.18958219606801116   0.6891295951078579   0.15927183297362668   0.4195989127928264   0.12666298206249849   0.24019508716665358   0.1400641193946152   0.8488914441986308   0.251630156674604   0.374006552248931   0.8570037322157779   0.9726164612735587   0.0011452616160246675
0.6395477491578472   0.8070509638423644   0.907799212263856   0.3508341703561695   0.5787622147544846   0.391976958510764   0.4887566578425655   0.45499875934541256   0.34602000170190494   0.1787572597953784   0.28777486329998897   0.2654165632774014   0.6568904065940471   0.019485426821751712   0.8681759505071626   0.1387535812149029   0.4166953194273935   0.8794213074271365   0.019284506308531797   0.8871234245402989   0.04268876717846252   0.022417575211358648   0.0466680450349731   0.8859781629242742   0.4031410180206153   0.2153666113689942   0.13886883277111717   0.5351439925681047   0.8243788032661307   0.8233896528582303   0.6501121749285517   0.08014523322269224   0.4783588015642258   0.6446323930628519   0.3623373116285627   0.8147286699452908   0.8214683949701787   0.6251469662411001   0.4941613611214001   0.6759750887303879   0.4047730755427852   0.7457256588139636   0.4748768548128683   0.788851664190089   0.36208430836432265   0.723308083602605   0.4282088097778952   0.9028735012658148   0.9589432903437074   0.5079414722336107   0.28933997700677805   0.36772950869771   0.13456448707757668   0.6845518193753806   0.6392278020782264   0.28758427547501775   0.6562056855133509   0.03991942631252864   0.2768904904496637   0.4728556055297269   0.8347372905431723   0.4147724600714285   0.7827291293282636   0.7968805167993389
0.42996421500038706   0.6690468012574649   0.3078522745153953   0.008028852609249935   0.06787990663606439   0.9457387176548598   0.8796434647375001   0.10515535134343518   0.10893661629235704   0.4377972454212491   0.590303487730722   0.7374258426457252   0.9743721292147803   0.7532454260458686   0.9510756856524957   0.44984156717070745   0.31816644370142944   0.71332599973334   0.674185195202832   0.9769859616409805   0.4834291531582572   0.29855353966191145   0.8914560658745685   0.18010544484164157   0.05346493815787012   0.6295067384044466   0.5836037913591732   0.17207659223239163   0.9855850315218058   0.6837680207495868   0.7039603266216731   0.06692124088895647   0.8766484152294487   0.2459707753283376   0.11365683889095099   0.32949539824323126   0.9022762860146684   0.492725349282469   0.1625811532384553   0.8796538310725238   0.5841098423132389   0.779399349549129   0.48839595803562325   0.9026678694315433   0.10068068915498174   0.4808458098872176   0.5969398921610548   0.7225624245899017   0.04721575099711161   0.851339071482771   0.013336100801881627   0.5504858323575101   0.06163071947530587   0.1675710507331843   0.30937577418020856   0.48356459146855363   0.18498230424585718   0.9216002754048467   0.19571893528925757   0.15406919322532234   0.28270601823118885   0.42887492612237765   0.033137782050802304   0.2744153621527985
0.6985961759179499   0.6494755765732485   0.5447418240151791   0.3717474927212552   0.5979154867629681   0.16862976668603094   0.9478019318541243   0.6491850681313535   0.5506997357658566   0.3172906952032599   0.9344658310522427   0.09869923577384337   0.4890690162905507   0.14971964447007563   0.6250900568720341   0.6151346443052897   0.3040867120446935   0.22811936906522898   0.4293711215827765   0.46106545107996744   0.021380693813504693   0.7992444429428514   0.3962333395319742   0.18665008892716892   0.3227845178955548   0.14976886636960282   0.8514915155167951   0.8149025962059138   0.7248690311325866   0.9811390996835719   0.9036895836626708   0.16571752807456025   0.17416929536673   0.663848404480312   0.9692237526104281   0.06701829230071689   0.6851002790761793   0.5141287600102363   0.3441336957383941   0.45188364799542713   0.3810135670314858   0.2860093909450073   0.9147625741556176   0.9908181969154597   0.3596328732179811   0.486764948002156   0.5185292346236434   0.8041681079882909   0.03684835532242633   0.3369960816325532   0.6670377191068483   0.9892655117823771   0.31197932418983976   0.35585698194898124   0.7633481354441775   0.8235479837078168   0.13781002882310972   0.6920085774686693   0.7941243828337492   0.7565296914070999   0.4527097497469304   0.17787981745843298   0.4499906870953551   0.3046460434116728
0.0716961827154446   0.8918704265134256   0.5352281129397375   0.3138278464962131   0.7120633094974635   0.40510547851126966   0.016698878316094116   0.5096597385079222   0.6752149541750372   0.06810939687871653   0.34966115920924584   0.5203942267255451   0.36323562998519743   0.7122524149297352   0.5863130237650684   0.6968462430177284   0.22542560116208774   0.020243837461065953   0.7921886409313191   0.9403165516106284   0.7727158514151573   0.842364020002633   0.342197953835964   0.6356705081989555   0.7010196686997127   0.9504935934892074   0.8069698408962265   0.3218426617027425   0.9889563592022492   0.5453881149779376   0.7902709625801324   0.8121829231948202   0.31374140502721204   0.4772787180992211   0.4406098033708865   0.29178869646927513   0.9505057750420146   0.7650263031694858   0.8542967796058182   0.5949424534515467   0.7250801738799268   0.7447824657084199   0.06210813867449899   0.6546259018409184   0.9523643224647695   0.9024184457057869   0.719910184838535   0.01895539364196281   0.2513446537650568   0.9519248522165796   0.9129403439423085   0.6971127319392203   0.2623882945628076   0.406536737238642   0.12266938136217612   0.8849298087444001   0.9486468895355956   0.9292580191394209   0.6820595779912896   0.5931411122751249   0.998141114493581   0.16423171596993502   0.8277627983854714   0.9981986588235782
0.27306094061365416   0.41944925026151514   0.7656546597109725   0.34357275698265977   0.3206966181488846   0.5170308045557283   0.04574447487243748   0.32461736334069696   0.06935196438382776   0.5651059523391486   0.132804130930129   0.6275046314014766   0.8069636698210202   0.15856921510050664   0.010134749567952869   0.7425748226570766   0.8583167802854246   0.22931119596108576   0.32807517157666327   0.1494337103819517   0.8601756657918436   0.06507947999115074   0.5003123731911918   0.15123505155837355   0.5871147251781894   0.6456302297296356   0.7346577134802194   0.8076622945757138   0.26641810702930485   0.12859942517390738   0.688913238607782   0.48304493123501685   0.1970661426454771   0.5634934728347588   0.556109107677653   0.8555402998335402   0.3901024728244569   0.4049242577342521   0.5459743581097001   0.11296547717646362   0.5317856925390324   0.17561306177316635   0.21789918653303678   0.9635317667945119   0.6716100267471887   0.11053358178201562   0.7175868133418449   0.8122967152361383   0.08449530156899934   0.46490335205238004   0.9829290998616256   0.004634420660424562   0.8180771945396945   0.33630392687847266   0.2940158612538436   0.5215894894254077   0.6210110518942175   0.7728104540437138   0.7379067535761906   0.6660491895918674   0.2309085790697605   0.3678861963094618   0.1919323954664906   0.5530837124154039
0.6991228865307282   0.1922731345362954   0.9740332089334538   0.589551945620892   0.02751285978353937   0.08173955275427978   0.2564463955916089   0.7772552303847535   0.94301755821454   0.6168362007018997   0.27351729572998335   0.772620809724329   0.12494036367484554   0.2805322738234271   0.9795014344761398   0.25103132029892133   0.5039293117806282   0.5077218197797132   0.24159468089994907   0.5849821307070538   0.27302073271086763   0.13983562347025144   0.049662285433458464   0.031898418291649994   0.5738978461801395   0.947562488933956   0.07562907650000464   0.44234647267075805   0.5463849863966   0.8658229361796762   0.8191826809083957   0.6650912422860045   0.60336742818206   0.2489867354777765   0.5456653851784123   0.8924704325616755   0.47842706450721456   0.9684544616543493   0.5661639507022727   0.6414391122627542   0.9744977527265865   0.4607326418746362   0.32456926980232353   0.05645698155570031   0.7014770200157188   0.3208970184043847   0.27490698436886507   0.02455856326405032   0.12757917383557935   0.37333452947042867   0.19927790786886043   0.5822120905932923   0.5811941874389792   0.5075115932907525   0.3800952269604647   0.9171208483072878   0.9778267592569192   0.2585248578129759   0.8344298417820524   0.024650415745612303   0.49939969474970464   0.2900703961586265   0.2682658910797797   0.38321130348285815
0.5249019420231182   0.8293377542839904   0.9436966212774561   0.3267543219271578   0.8234249220073994   0.5084407358796057   0.6687896369085911   0.3021957586631075   0.6958457481718201   0.13510620640917698   0.46951172903973065   0.7199836680698153   0.11465156073284084   0.6275946131184246   0.08941650207926595   0.8028628197625275   0.1368248014759217   0.3690697553054486   0.2549866602972136   0.7782124040169152   0.637425106726217   0.07899935914682209   0.9867207692174339   0.395001100534057   0.11252316470309884   0.24966160486283173   0.04302414793997771   0.06824677860689919   0.28909824269569945   0.741220868983226   0.3742345110313866   0.7660510199437917   0.5932524945238794   0.6061146625740491   0.9047227819916559   0.046067351873976425   0.4786009337910385   0.9785200494556245   0.81530627991239   0.24320453211144896   0.34177613231511683   0.6094502941501759   0.5603196196151764   0.4649921280945338   0.7043510255888998   0.5304509350033538   0.5735988503977425   0.06999102756047675   0.591827860885801   0.2807893301405221   0.5305747024577647   0.0017442489535775519   0.3027296181901015   0.5395684611572961   0.15634019142637817   0.23569322900978587   0.7094771236662222   0.933453798583247   0.2516174094347222   0.18962587713580945   0.23087618987518363   0.9549337491276224   0.43631112952233225   0.9464213450243605
0.8891000575600668   0.3454834549774464   0.8759915099071559   0.4814292169298267   0.184749031971167   0.8150325199740927   0.30239265950941335   0.41143818936934995   0.592921171085366   0.5342431898335704   0.7718179570516486   0.40969394041577245   0.2901915528952645   0.9946747286762745   0.6154777656252705   0.17400071140598655   0.5807144292290424   0.06122093009302751   0.3638603561905482   0.9843748342701771   0.3498382393538587   0.10628718096540514   0.9275492266682159   0.0379534892458166   0.46073818179379195   0.7608037259879586   0.05155771676106011   0.5565242723159899   0.27598914982262496   0.9457712060138661   0.7491650572516467   0.1450860829466399   0.6830679787372589   0.4115280161802956   0.9773471001999982   0.7353921425308675   0.3928764258419944   0.4168532875040212   0.3618693345747277   0.5613914311248809   0.8121619966129521   0.3556323574109937   0.9980089783841795   0.5770165968547039   0.4623237572590933   0.24934517644558854   0.07045975171596353   0.5390631076088872   0.0015855754653013782   0.48854145045762987   0.01890203495490342   0.9825388352928973   0.7255964256426765   0.5427702444437638   0.26973697770325666   0.8374527523462575   0.04252844690541754   0.13124222826346812   0.29238987750325857   0.10206060981538996   0.6496520210634231   0.7143889407594469   0.9305205429285308   0.540669178690509
0.8374900244504712   0.3587565833484533   0.9325115645443514   0.9636525818358052   0.3751662671913778   0.10941140690286474   0.8620518128283878   0.42458947422691795   0.37358069172607644   0.6208699564452349   0.8431497778734844   0.44205063893402063   0.6479842660834   0.07809971200147114   0.5734128001702278   0.6045978865877631   0.6054558191779824   0.946857483738003   0.28102292266696915   0.5025372767723733   0.9558037981145593   0.23246854297855607   0.3505023797384383   0.9618680980818642   0.1183137736640882   0.8737119596301027   0.41799081519408693   0.998215516246059   0.7431475064727104   0.7643005527272381   0.555939002365699   0.573626042019141   0.36956681474663394   0.14343059628200314   0.7127892244922147   0.1315754030851204   0.721582548663234   0.06533088428053198   0.13937642432198694   0.5269775164973572   0.11612672948525153   0.11847340054252897   0.8583535016550178   0.024440239724983992   0.16032293137069223   0.886004857563973   0.5078511219165794   0.06257214164311979   0.04200915770660403   0.012292897933870138   0.0898603067224925   0.06435662539706079   0.29886165123389363   0.2479923452066321   0.5339213043567934   0.49073058337791975   0.9292948364872596   0.10456174892462898   0.8211320798645787   0.35915518029279936   0.2077122878240257   0.03923086464409699   0.6817556555425918   0.8321776637954421
0.09158555833877416   0.920757464101568   0.8234021538875741   0.8077374240704581   0.9312626269680819   0.034752606537595106   0.3155510319709946   0.7451652824273384   0.8892534692614779   0.022459708603724968   0.22569072524850212   0.6808086570302776   0.5903918180275842   0.7744673633970929   0.6917694208917087   0.1900780736523578   0.6610969815403246   0.6699056144724639   0.87063734102713   0.8309228933595584   0.4533846937162989   0.6306747498283669   0.18888168548453815   0.9987452295641163   0.3617991353775247   0.7099172857267989   0.3654795315969641   0.19100780549365814   0.4305365084094428   0.6751646791892038   0.04992849962596949   0.4458425230663198   0.5412830391479649   0.6527049705854788   0.8242377743774674   0.7650338660360423   0.9508912211203806   0.878237607188386   0.1324683534857587   0.5749557923836844   0.289794239580056   0.20833199271592207   0.2618310124586287   0.7440328990241261   0.8364095458637572   0.5776572428875552   0.07294932697409058   0.7452876694600097   0.47461041048623237   0.8677399571607562   0.7074697953771265   0.5542798639663515   0.04407390207678956   0.19257527797155252   0.6575412957511569   0.10843734090003178   0.5027908629288247   0.5398703073860738   0.8333035213736896   0.34340347486398953   0.5518996418084441   0.6616327001976878   0.7008351678879309   0.768447682480305
0.262105402228388   0.4533007074817657   0.43900415542930216   0.024414783456179076   0.4256958563646309   0.8756434645942106   0.3660548284552116   0.27912711399616935   0.9510854458783986   0.00790350743345427   0.6585850330780851   0.7248472500298178   0.907011543801609   0.8153282294619018   0.0010437373269281285   0.616409909129786   0.40422068087278434   0.27545792207582803   0.16774021595323851   0.27300643426579646   0.8523210390643403   0.6138252218781403   0.46690504806530764   0.5045587517854914   0.5902156368359522   0.1605245143963745   0.027900892636005425   0.48014396832931233   0.16451978047132135   0.28488104980216394   0.6618460641807938   0.20101685433314295   0.2134343345929228   0.27697754236870964   0.0032610311027087054   0.47616960430332517   0.3064227907913138   0.4616493129068079   0.0022172937757805765   0.8597596951735391   0.9022021099185294   0.1861913908309799   0.8344770778225421   0.5867532609077427   0.04988107085418919   0.5723661689528396   0.36757202975723446   0.08219450912225128   0.45966543401823695   0.4118416545564652   0.33967113712122904   0.602050540792939   0.2951456535469156   0.12696060475430127   0.6778250729404351   0.401033686459796   0.08171131895399279   0.8499830623855916   0.6745640418377264   0.9248640821564709   0.775288528162679   0.3883337494787837   0.6723467480619459   0.06510438698293167
0.8730864182441496   0.2021423586478038   0.8378696702394038   0.478351126075189   0.8232053473899603   0.6297761896949641   0.47029764048216943   0.3961566169529377   0.36353991337172337   0.21793453513849892   0.1306265033609404   0.7941060761599987   0.0683942598248078   0.09097393038419767   0.4528014304205052   0.39307238970020275   0.986682940870815   0.24099086799860606   0.7782373885827787   0.46820830754373194   0.21139441270813603   0.8526571185198224   0.10589064052083282   0.40310392056080024   0.3383079944639865   0.6505147598720186   0.26802097028142896   0.9247527944856113   0.5151026470740262   0.020738570177054418   0.7977233297992595   0.5285961775326735   0.15156273370230278   0.8028040350385555   0.6670968264383191   0.7344901013726748   0.08316847387749497   0.7118301046543578   0.21429539601781394   0.3414177116724721   0.09648553300667997   0.4708392366557518   0.4360580074350352   0.8732094041287402   0.885091120298544   0.6181821181359294   0.3301673669142024   0.4701054835679399   0.5467831258345575   0.9676673582639109   0.062146396632773444   0.5453526890823286   0.031680478760531275   0.9469287880868564   0.2644230668335139   0.016756511549655073   0.8801177450582285   0.144124753048301   0.5973262403951948   0.28226641017698023   0.7969492711807336   0.43229464839394316   0.38303084437738083   0.9408486985045081
0.7004637381740535   0.9614554117381914   0.9469728369423456   0.06763929437576797   0.8153726178755096   0.34327329360226194   0.6168054700281432   0.5975338108078281   0.26858949204095217   0.37560593533835107   0.5546590733953698   0.05218112172549942   0.23690901328042088   0.4286771472514946   0.29023600656185583   0.03542461017584435   0.35679126822219237   0.2845523942031936   0.6929097661666611   0.7531581999988641   0.5598419970414589   0.8522577458092505   0.3098789217892803   0.812309501494356   0.8593782588674054   0.890802334071059   0.36290608484693465   0.744670207118588   0.04400564099189574   0.5475290404687971   0.7461006148187914   0.14713639631075992   0.7754161489509436   0.17192310513044604   0.19144154142342173   0.0949552745852605   0.5385071356705227   0.7432459578789514   0.9012055348615658   0.059530664409416144   0.18171586744833032   0.4586935636757578   0.2082957686949048   0.30637246441055205   0.6218738704068715   0.6064358178665074   0.8984168469056245   0.49406296291619606   0.7624956115394661   0.7156334837954482   0.5355107620586899   0.7493927557976081   0.7184899705475704   0.16810444332665114   0.7894101472398983   0.6022563594868482   0.9430738215966268   0.9961813381962051   0.5979686058164766   0.5073010849015877   0.40456668592610406   0.2529353803172537   0.6967630709549107   0.44777042049217153
0.22285081847777374   0.7942418166414958   0.488467302260006   0.1413979560816195   0.6009769480709023   0.18780599877498855   0.5900504553543815   0.6473349931654234   0.8384813365314362   0.47217251497954027   0.05453969329569163   0.8979422373678153   0.1199913659838658   0.3040680716528891   0.26512954605579325   0.2956858778809672   0.176917544387239   0.30788673345668405   0.6671609402393166   0.7883847929793795   0.7723508584611349   0.05495135313943033   0.9703978692844059   0.34061437248720794   0.5495000399833612   0.26070953649793444   0.4819305670243999   0.19921641640558843   0.9485230919124589   0.07290353772294589   0.8918801116700183   0.551881423240165   0.11004175538102268   0.6007310227434056   0.8373404183743268   0.6539391858723497   0.9900503893971568   0.29666295109051644   0.5722108723185335   0.3582533079913825   0.8131328450099179   0.9887762176338324   0.9050499320792169   0.569868515012003   0.04078198654878297   0.933824864494402   0.9346520627948111   0.22925414252479503   0.4912819465654218   0.6731153279964677   0.45272149577041115   0.03003772611920662   0.5427588546529629   0.6002117902735218   0.5608413841003927   0.47815630287904165   0.4327170992719403   0.9994807675301162   0.7235009657260659   0.824217117006692   0.4426667098747834   0.7028178164395997   0.15129009340753247   0.46596380901530954
0.6295338648648655   0.7140415988057673   0.24624016132831558   0.8960952940033066   0.5887518783160826   0.7802167343113652   0.31158809853350455   0.6668411514785115   0.09746993175066072   0.10710140631489755   0.8588666027630935   0.6368034253593049   0.5547110770976977   0.5068896160413757   0.29802521866270065   0.15864712248026325   0.1219939778257575   0.5074088485112596   0.5745242529366347   0.33443000547357127   0.6793272679509741   0.8045910320716598   0.42323415952910226   0.8684661964582617   0.04979340308610859   0.09054943326589256   0.17699399820078665   0.9723709024549552   0.4610415247700261   0.31033269895452736   0.8654058996672821   0.3055297509764437   0.3635715930193653   0.2032312926396298   0.006539296904188684   0.6687263256171389   0.8088605159216675   0.6963416765982541   0.708514078241488   0.5100792031368756   0.68686653809591   0.18893282808699444   0.13398982530485332   0.17564919766330434   0.007539270144935965   0.3843417960153346   0.7107556657757511   0.3071830012050426   0.9577458670588274   0.29379236274944204   0.5337616675749643   0.33481209875008744   0.49670434228880134   0.9834596637949147   0.6683557679076823   0.029282347773643753   0.133132749269436   0.7802283711552849   0.6618164710034936   0.36055602215650495   0.32427223334776845   0.08388669455703085   0.9533023927620056   0.8504768190196293
0.6374056952518584   0.8949538664700364   0.8193125674571523   0.674827621356325   0.6298664251069224   0.5106120704547018   0.10855690168140124   0.36764462015128235   0.672120558048095   0.21681970770525982   0.5747952341064368   0.03283252140119492   0.1754162157592937   0.23336004391034515   0.9064394661987545   0.0035501736275511658   0.042283466489857716   0.4531316727550603   0.24462299519526093   0.6429941514710462   0.7180112331420893   0.3692449781980294   0.2913206024332553   0.7925173324514169   0.08060553789023091   0.474291111727993   0.472008034976103   0.1176897110950919   0.45073911278330847   0.9636790412732912   0.36345113329470174   0.7500450909438096   0.7786185547352135   0.7468593335680314   0.788655899188265   0.7172125695426146   0.6032023389759198   0.5134992896576862   0.8822164329895104   0.7136623959150634   0.560918872486062   0.06036761690262593   0.6375934377942495   0.0706682444440172   0.8429076393439727   0.6911226387045966   0.3462728353609942   0.27815091199260034   0.7623021014537419   0.21683152697660352   0.8742648003848912   0.16046120089750843   0.31156298867043336   0.25315248570331234   0.5108136670901894   0.41041610995369887   0.53294443393522   0.506293152135281   0.7221577679019244   0.6932035404110843   0.9297420949593002   0.9927938624775948   0.8399413349124141   0.9795411444960208
0.3688232224732381   0.9324262455749689   0.2023478971181646   0.9088729000520036   0.5259155831292653   0.24130360687037236   0.8560750617571704   0.6307219880594034   0.7636134816755235   0.024472079893768855   0.9818102613722792   0.4702607871618949   0.45205049300509015   0.7713195941904565   0.4709965942820899   0.05984467720819603   0.9191060590698702   0.2650264420551755   0.7488388263801654   0.36664113679711174   0.98936396411057   0.2722325795775807   0.9088974914677513   0.3870999923010909   0.620540741637332   0.33980633400261184   0.7065495943495868   0.4782270922490872   0.09462515850806663   0.09850272713223945   0.8504745325924163   0.8475051041896838   0.3310116768325431   0.07403064723847061   0.8686642712201371   0.37724431702778893   0.878961183827453   0.3027110530480141   0.3976676769380472   0.3173996398195929   0.9598551247575827   0.037684610992838596   0.6488288505578818   0.9507585030224812   0.9704911606470127   0.7654520314152579   0.7399313590901304   0.5636585107213903   0.34995041900968066   0.4256456974126461   0.033381764740543586   0.08543141847230308   0.255325260501614   0.3271429702804066   0.1829072321481272   0.2379263142826192   0.9243135836690709   0.25311232304193604   0.3142429609279901   0.8606819972548303   0.04535239984161793   0.9504012699939219   0.9165752839899429   0.5432823574352373
0.08549727508403518   0.9127166590010833   0.2677464334320611   0.5925238544127561   0.11500611443702252   0.14726462758582543   0.5278150743419308   0.028865343691365845   0.7650556954273419   0.7216189301731794   0.4944333096013871   0.9434339252190628   0.5097304349257278   0.39447595989277273   0.31152607745325994   0.7055076109364435   0.5854168512566569   0.1413636368508367   0.9972831165252698   0.8448256136816132   0.5400644514150389   0.19096236685691476   0.08070783253532694   0.30154325624637596   0.45456717633100374   0.2782457078558314   0.8129613991032658   0.7090194018336198   0.3395610618939812   0.13098108027000602   0.2851463247613351   0.6801540581422539   0.5745053664666394   0.40936215009682664   0.790713015159948   0.7367201329231912   0.0647749315409116   0.014886190204053944   0.4791869377066881   0.031212521986747645   0.47935808028425475   0.8735225533532173   0.4819038211814183   0.18638690830513435   0.9392936288692159   0.6825601864963025   0.40119598864609135   0.8848436520587584   0.48472645253821206   0.40431447864047104   0.5882345895428255   0.17582425022513862   0.14516539064423084   0.27333339837046505   0.30308826478149037   0.49567019208288465   0.5706600241775914   0.8639712482736384   0.5123752496215424   0.7589500591596935   0.5058850926366798   0.8490850580695845   0.033188311914854246   0.7277375371729459
0.026527012352425088   0.9755625047163672   0.551284490733436   0.5413506288678115   0.08723338348320928   0.2930023182200647   0.15008850208734462   0.656506976809053   0.6025069309449972   0.8886878395795936   0.5618539125445191   0.4806827265839144   0.45734154030076635   0.6153544412091286   0.2587656477630288   0.9850125345010298   0.8866815161231749   0.7513831929354903   0.7463903981414864   0.2260624753413363   0.3807964234864951   0.9022981348659058   0.7132020862266322   0.49832493816839046   0.35426941113407   0.9267356301495386   0.1619175954931962   0.956974309300579   0.2670360276508607   0.6337333119294739   0.011829093405851594   0.3004673324915259   0.6645290967058636   0.7450454723498803   0.4499751808613325   0.8197846059076115   0.20718755640509715   0.12969103114075167   0.1912095330983037   0.8347720714065817   0.3205060402819222   0.3783078382052614   0.4448191349568173   0.6087095960652454   0.9397096167954271   0.4760097033393556   0.7316170487301851   0.11038465789685493   0.5854402056613571   0.5492740731898169   0.5696994532369889   0.15341034859627595   0.3184041780104964   0.915540761260343   0.5578703598311373   0.85294301610475   0.6538750813046329   0.17049528891046267   0.10789517896980481   0.033158410197138534   0.4466875248995357   0.040804257769711   0.9166856458715011   0.19838633879055684
0.1261814846176135   0.6624964195644496   0.47186651091468385   0.5896767427253115   0.18647186782218636   0.18648671622509397   0.7402494621844987   0.4792920848284565   0.6010316621608293   0.637212643035277   0.17055000894750985   0.32588173623218053   0.28262748415033284   0.721671881774934   0.6126796491163726   0.4729387201274305   0.6287524028457   0.5511765928644713   0.5047844701465678   0.439780309930292   0.18206487794616424   0.5103723350947603   0.5880988242750667   0.24139397113973515   0.05588339332855074   0.8478759155303107   0.1162323133603828   0.6517172284144237   0.8694115255063644   0.6613891993052168   0.37598285117588404   0.17242514358596725   0.26837986334553515   0.024176556269939777   0.20543284222837419   0.8465434073537867   0.9857523791952023   0.30250467449500573   0.5927531931120016   0.3736046872263562   0.35699997634950237   0.7513280816305344   0.08796872296543386   0.9338243772960643   0.17493509840333815   0.24095574653577406   0.49986989869036724   0.6924304061563291   0.1190517050747874   0.3930798310054633   0.38363758532998443   0.040713177741905346   0.24964017956842302   0.7316906317002465   0.00765473415410038   0.8682880341559381   0.9812603162228879   0.7075140754303068   0.8022218919257262   0.02174462680215136   0.9955079370276855   0.40500940093530097   0.20946869881372457   0.6481399395757952
0.6385079606781832   0.6536813193047666   0.12149997584829071   0.7143155622797309   0.463572862274845   0.4127255727689925   0.6216300771579235   0.021885156123401833   0.3445211572000576   0.019645741763529227   0.23799249182793905   0.9811719783814965   0.0948809776316346   0.2879551100632827   0.23033775767383868   0.1128839442255584   0.11362066140874673   0.580441034632976   0.4281158657481125   0.09113931742340704   0.1181127243810612   0.17543163369767506   0.2186471669343879   0.4429993778476119   0.4796047637028781   0.5217503143929085   0.09714719108609719   0.728683815567881   0.01603190142803304   0.10902474162391597   0.4755171139281737   0.7067986594444792   0.6715107442279754   0.08937899986038675   0.23752462210023467   0.7256266810629827   0.5766297665963408   0.801423889797104   0.007186864426395993   0.6127427368374243   0.4630091051875941   0.22098285516412797   0.5790709986782835   0.5216034194140172   0.3448963808065329   0.04555122146645292   0.3604238317438956   0.07860404156640531   0.8652916171036549   0.5238009070735444   0.2632766406577984   0.3499202259985243   0.8492597156756219   0.4147761654496285   0.7877595267296247   0.6431215665540452   0.17774897144764637   0.3253971655892417   0.5502349046293901   0.9174948854910625   0.6011192048513055   0.5239732757921377   0.543048040202994   0.30475214865363826
0.13811009966371143   0.30299042062800974   0.9639770415247105   0.783148729239621   0.7932137188571785   0.25743919916155683   0.603553209780815   0.7045446876732157   0.9279221017535236   0.7336382920880123   0.3402765691230165   0.35462446167469136   0.07866238607790187   0.3188621266383839   0.5525170423933918   0.7115028951206462   0.9009134146302555   0.9934649610491422   0.0022821377640018068   0.7940080096295837   0.29979420977894994   0.46949168525700447   0.4592340975610078   0.4892558609759455   0.16168411011523853   0.16650126462899476   0.49525705603629727   0.7061071317363244   0.36847039125806   0.909062065467438   0.8917038462554824   0.0015624440631087841   0.44054828950453634   0.17542377337942558   0.5514272771324659   0.6469379823884174   0.36188590342663446   0.8565616467410416   0.998910234739074   0.9354350872677711   0.460972488796379   0.8630966856918995   0.9966280969750722   0.14142707763818746   0.161178279017429   0.393605000434895   0.5373939994140644   0.652171216662242   0.9994941689021904   0.22710373580590024   0.042136943377767154   0.9460640849259174   0.6310237776441304   0.3180416703384623   0.1504330971222848   0.9445016408628086   0.19047548813959414   0.14261789695903673   0.5990058199898189   0.29756365847439126   0.8285895847129596   0.2860562502179951   0.600095585250745   0.3621285712066201
0.3676170959165807   0.42295956452609557   0.6034674882756728   0.22070149356843266   0.2064388168991517   0.029354564091200578   0.0660734888616084   0.5685302769061907   0.20694464799696122   0.8022508282853004   0.023936545483841234   0.6224661919802732   0.5759208703528307   0.48420915794683805   0.8735034483615565   0.6779645511174646   0.3854453822132366   0.3415912609878013   0.2744976283717374   0.3804008926430733   0.5568557975002769   0.05553501076980625   0.6744020431209925   0.018272321436453194   0.1892387015836962   0.6325754462437106   0.07093455484531964   0.7975708278680206   0.9827998846845445   0.6032208821525101   0.004861065983711256   0.22904055096182985   0.7758552366875833   0.8009700538672098   0.98092452049987   0.6065743589815566   0.1999343663347526   0.3167608959203717   0.10742107213831359   0.9286098078640921   0.814488984121516   0.9751696349325705   0.8329234437665761   0.5482089152210188   0.2576331866212391   0.9196346241627642   0.1585214006455837   0.5299365937845656   0.06839448503754286   0.2870591779190535   0.08758684580026406   0.732365765916545   0.08559460035299835   0.6838382957665434   0.08272577981655281   0.5033252149547152   0.30973936366541505   0.8828682418993337   0.10180125931668278   0.8967508559731585   0.10980499733066244   0.566107345978962   0.9943801871783692   0.9681410481090665
0.29531601320914647   0.5909377110463915   0.16145674341179303   0.41993213288804776   0.037682826587907364   0.6713030868836273   0.002935342766209325   0.8899955391034822   0.9692883415503645   0.38424390896457383   0.9153484969659452   0.1576297731869372   0.8836937411973662   0.7004056131980304   0.8326227171493924   0.654304558232222   0.5739543775319511   0.8175373712986967   0.7308214578327097   0.7575537022590635   0.4641493802012887   0.25143002531973485   0.7364412706543405   0.789412654149997   0.16883336699214224   0.6604923142733433   0.5749845272425474   0.3694805212619492   0.13115054040423488   0.989189227389716   0.5720491844763381   0.479484982158467   0.16186219885387038   0.6049453184251422   0.6567006875103929   0.3218552089715298   0.2781684576565042   0.9045397052271118   0.8240779703610004   0.6675506507393077   0.7042140801245531   0.08700233392841504   0.09325651252829073   0.9099969484802443   0.2400646999232644   0.8355723086086801   0.35681524187395025   0.12058429433024731   0.07123133293112215   0.17507999433533686   0.7818307146314029   0.7511037730682981   0.9400807925268873   0.18589076694562082   0.20978153015506473   0.2716187909098311   0.7782185936730169   0.5809454485204786   0.5530808426446718   0.9497635819383013   0.5000501360165127   0.6764057432933668   0.7290028722836714   0.28221293119899354
0.7958360558919596   0.5894034093649517   0.6357463597553807   0.3722159827187493   0.5557713559686952   0.7538311007562716   0.2789311178814305   0.251631688388502   0.48454002303757304   0.5787511064209347   0.49710040325002763   0.5005279153202039   0.5444592305106858   0.3928603394753139   0.2873188730949629   0.22890912441037278   0.7662406368376689   0.8119148909548353   0.734238030450291   0.27914554247207146   0.2661905008211562   0.1355091476614685   0.005235158166619556   0.996932611273078   0.47035444492919665   0.5461057382965168   0.36948879841123883   0.6247166285543286   0.9145830889605014   0.7922746375402452   0.09055768052980832   0.37308494016582666   0.43004306592292846   0.21352353111931047   0.5934572772797807   0.8725570248456228   0.8855838354122427   0.8206631916439966   0.30613840418481775   0.64364790043525   0.11934319857457384   0.008748300689161263   0.5719003737345267   0.3645023579631786   0.8531526977534176   0.8732391530276927   0.5666652155679072   0.3675697466901007   0.38279825282422103   0.327133414731176   0.19717641715666837   0.742853118135772   0.46821516386371953   0.5348587771909309   0.10661873662686003   0.3697681779699453   0.038172097940791086   0.3213352460716204   0.5131614593470794   0.4972111531243225   0.15258826252854837   0.5006720544276239   0.2070230551622616   0.8535632526890725
0.03324506395397454   0.4919237537384626   0.6351226814277349   0.4890608947258939   0.1800923662005569   0.6186846007107698   0.0684574658598277   0.12149114803579325   0.7972941133763359   0.2915511859795938   0.8712810487031594   0.37863802990002127   0.32907894951261635   0.756692408788663   0.7646623120762993   0.008869851930075917   0.2909068515718253   0.43535716271704256   0.25150085272921996   0.5116586988057534   0.1383185890432769   0.9346851082894188   0.044477797566958376   0.6580954461166809   0.10507352508930236   0.4427613545509561   0.4093551161392235   0.16903455139078702   0.9249811588887454   0.8240767538401863   0.3408976502793958   0.047543403354993755   0.12768704551240956   0.5325255678605926   0.4696166015762364   0.6689053734549725   0.7986080959997932   0.7758331590719296   0.7049542894999371   0.6600355215248966   0.5077012444279679   0.3404759963548871   0.45345343677071714   0.14837682271914318   0.369382655384691   0.40579088806546837   0.4089756392037588   0.4902813766024623   0.26430913029538866   0.9630295335145123   0.9996205230645353   0.32124682521167525   0.3393279714066432   0.13895277967432593   0.6587228727851395   0.2737034218566815   0.21164092589423364   0.6064272118137334   0.18910627120890305   0.604798048401709   0.41303282989444046   0.8305940527418038   0.48415198170896595   0.9447625268768124
0.9053315854664725   0.49011805638691663   0.03069854493824877   0.7963857041576692   0.5359489300817815   0.08432716832144824   0.62172290573449   0.30610432755520695   0.2716397997863928   0.12129763480693599   0.6221023826699548   0.9848575023435316   0.9323118283797496   0.98234485513261   0.9633795098848152   0.7111540804868501   0.7206709024855159   0.3759176433188767   0.7742732386759121   0.10635603208514115   0.3076380725910755   0.545323590577073   0.29012125696694624   0.1615935052083287   0.40230648712460304   0.055205534190156336   0.2594227120286975   0.3652078010506595   0.8663575570428216   0.9708783658687081   0.6376998062942075   0.05910347349545254   0.5947177572564287   0.8495807310617721   0.015597423624252784   0.07424597115192086   0.6624059288766792   0.8672358759291621   0.05221791373943755   0.3630918906650707   0.9417350263911631   0.49131823261028534   0.2779446750635254   0.25673585857992953   0.6340969538000877   0.9459946420332124   0.9878234180965791   0.09514235337160083   0.2317904666754846   0.890789107843056   0.7284007060678817   0.7299345523209413   0.3654329096326631   0.919910741974348   0.09070089977367411   0.6708310788254888   0.7707151523762343   0.07033001091257582   0.07510347614942132   0.596585107673568   0.10830922349955525   0.20309413498341378   0.022885562409983767   0.23349321700849723
0.16657419710839208   0.7117759023731285   0.7449408873464584   0.9767573584285677   0.5324772433083045   0.7657812603399161   0.7571174692498793   0.8816150050569669   0.30068677663281984   0.87499215249686   0.028716763181997694   0.1516804527360255   0.9352538670001568   0.9550814105225122   0.9380158634083235   0.4808493739105367   0.16453871462392236   0.8847513996099363   0.8629123872589023   0.8842642662369687   0.05622949112436713   0.6816572646265225   0.8400268248489184   0.6507710492284715   0.889655294015975   0.969881362253394   0.0950859375024601   0.6740136907999038   0.35717805070767056   0.204100101913478   0.3379684682525808   0.792398685742937   0.05649127407485075   0.3291079494166179   0.3092517050705831   0.6407182330069114   0.121237407074694   0.3740265388941058   0.37123584166225954   0.15986885909637474   0.9566986924507717   0.4892751392841695   0.5083234544033572   0.275604592859406   0.9004692013264045   0.8076178746576469   0.6682966295544388   0.6248335436309344   0.010813907310429475   0.8377365124042528   0.5732106920519786   0.9508198528310305   0.6536358566027589   0.6336364104907748   0.23524222379939785   0.15842116708809356   0.5971445825279081   0.3045284610741569   0.9259905187288148   0.5177029340811821   0.47590717545321415   0.9305019221800511   0.5547546770665552   0.35783407498480735
0.5192084830024425   0.44122678289588163   0.046431222663198005   0.08222948212540139   0.618739281676038   0.6336089082382347   0.37813459310875924   0.45739593849446697   0.6079253743656086   0.7958723958339818   0.8049239010567806   0.5065760856634365   0.9542895177628496   0.16223598534320707   0.5696816772573827   0.34815491857534286   0.35714493523494145   0.8577075242690502   0.643691158528568   0.8304519844941608   0.8812377597817274   0.9272056020889992   0.0889364814620127   0.47261790950935345   0.36202927677928487   0.4859788191931175   0.0425052587988147   0.3903884273839521   0.7432899951032469   0.8523699109548828   0.6643706656900554   0.932992488889485   0.13536462073763836   0.056497515120900905   0.8594467646332749   0.4264164032260486   0.18107510297478874   0.8942615297776938   0.2897650873758921   0.07826148465070575   0.8239301677398473   0.03655400550864365   0.6460739288473242   0.24780950015654496   0.9426924079581199   0.10934840341964454   0.5571374473853115   0.7751915906471916   0.5806631311788351   0.623369584226527   0.5146321885864967   0.38480316326323943   0.8373731360755882   0.7709996732716443   0.8502615228964413   0.4518106743737544   0.7020085153379498   0.7145021581507434   0.9908147582631665   0.02539427114770576   0.520933412363161   0.8202406283730496   0.7010496708872743   0.9471327864970001
0.6970032446233139   0.7836866228644058   0.05497574203995016   0.699323286340455   0.7543108366651939   0.6743382194447614   0.4978382946546387   0.9241316956932636   0.17364770548635883   0.05096863521823428   0.983206106068142   0.5393285324300241   0.33627456941077066   0.27996896194659004   0.1329445831717006   0.08751785805626969   0.6342660540728208   0.5654668037958467   0.14212982490853415   0.06212358690856393   0.11333264170965972   0.7452261754227971   0.44108015402125983   0.11499080041156391   0.41632939708634586   0.9615395525583913   0.3861044119813096   0.41566751407110886   0.662018560421152   0.28720133311362994   0.8882661173266709   0.4915358183778453   0.48837085493479315   0.23623269789539567   0.9050600112585291   0.9522072859478212   0.15209628552402252   0.9562637359488056   0.7721154280868284   0.8646894278915516   0.5178302314512017   0.39079693215295896   0.6299856031782943   0.8025658409829877   0.404497589741542   0.6455707567301618   0.18890544915703447   0.6875750405714237   0.9881681926551961   0.6840312041717705   0.8028010371757248   0.27190752650031486   0.32614963223404414   0.3968298710581406   0.9145349198490539   0.7803717081224695   0.837778777299251   0.1605971731627449   0.009474908590524824   0.8281644221746483   0.6856824917752284   0.20433343721393926   0.2373594805036964   0.9634749942830967
0.16785226032402675   0.8135365050609803   0.6073738773254022   0.1609091533001091   0.7633546705824847   0.16796574833081845   0.41846842816836766   0.4733341127286854   0.7751864779272887   0.4839345441590479   0.6156673909926429   0.20142658622837056   0.44903684569324454   0.08710467310090733   0.701132471143589   0.42105487810590103   0.6112580683939935   0.9265074999381624   0.6916575625530642   0.5928904559312528   0.9255755766187651   0.7221740627242231   0.4542980820493678   0.629415461648156   0.7577233162947383   0.9086375576632428   0.8469242047239657   0.4685063083480469   0.9943686457122536   0.7406718093324244   0.42845577655559797   0.9951721956193615   0.2191821677849649   0.25673726517337647   0.8127883855629552   0.7937456093909909   0.7701453220917204   0.16963259207246914   0.11165591441936615   0.3726907312850899   0.15888725369772683   0.24312509213430672   0.41999835186630197   0.7798002753538371   0.23331167707896172   0.5209510294100835   0.9657002698169342   0.1503848137056811   0.4755883607842234   0.6123134717468407   0.11877606509296859   0.6818785053576342   0.4812197150719698   0.8716416624144163   0.6903202885373706   0.6867063097382727   0.2620375472870049   0.6149043972410398   0.8775319029744155   0.8929607003472818   0.4918922251952845   0.4452718051685707   0.7658759885550493   0.5202699690621919
0.3330049714975577   0.202146713034264   0.3458776366887473   0.7404696937083548   0.09969329441859598   0.6811956836241805   0.3801773668718131   0.5900848800026737   0.6241049336343726   0.06888221187733973   0.2614013017788445   0.9082063746450394   0.1428852185624028   0.1972405494629234   0.5710810132414739   0.22150006490676674   0.880847671275398   0.5823361522218836   0.6935491102670585   0.32853936455948496   0.38895544608011345   0.13706434705331288   0.9276731217120091   0.808269395497293   0.05595047458255574   0.9349176340190489   0.5817954850232617   0.06779970178893834   0.9562571801639598   0.25372195039486845   0.20161811815144867   0.4777148217862647   0.33215224652958714   0.18483973851752875   0.9402168163726041   0.5695084471412253   0.18926702796718434   0.9875991890546053   0.3691358031311303   0.3480083822344585   0.30841935669178644   0.40526303683272175   0.6755866928640719   0.01946901767497353   0.919463910611673   0.26819868977940886   0.7479135711520628   0.21119962217768043   0.8635134360291172   0.33328105576036   0.16611808612880102   0.1433999203887421   0.9072562558651575   0.07955910536549152   0.9644999679773524   0.6656850986024774   0.5751040093355704   0.8947193668479628   0.024283151604748168   0.09617665146125216   0.385836981368386   0.9071201777933574   0.6551473484736179   0.7481682692267937
0.07741762467659957   0.5018571409606357   0.979560655609546   0.7286992515518201   0.1579537140649266   0.23365845118122686   0.23164708445748322   0.5174996293741397   0.2944402780358093   0.9003773954208669   0.0655289983286822   0.37409970898539757   0.38718402217065184   0.8208182900553753   0.10102903035132985   0.7084146103829202   0.8120800128350815   0.9260989232074126   0.07674587874658167   0.612237958921668   0.4262430314666955   0.01897874541405512   0.4215985302729638   0.8640696896948744   0.34882540679009594   0.5171216044534194   0.4420378746634178   0.13537043814305424   0.19087169272516935   0.28346315327219257   0.2103907902059346   0.6178708087689145   0.89643141468936   0.3830857578513257   0.1448617918772524   0.243771099783517   0.5092473925187082   0.5622674677959504   0.04383276152592255   0.5353564894005968   0.6971673796836267   0.6361685445885378   0.9670868827793409   0.9231185304789288   0.2709243482169312   0.6171897991744827   0.5454883525063771   0.05904884078405442   0.9220989414268352   0.10006819472106324   0.10345047784295927   0.9236784026410002   0.7312272487016659   0.8166050414488707   0.8930596876370247   0.3058075938720856   0.834795834012306   0.433519283597545   0.7481978957597722   0.06203649408856863   0.32554844149359774   0.8712518158015946   0.7043651342338497   0.5266800046879718
0.628381061809971   0.2350832712130569   0.7372782514545089   0.603561474209043   0.3574567135930398   0.6178934720385743   0.19178989894813178   0.5445126334249886   0.4353577721662045   0.517825277317511   0.0883394211051725   0.6208342307839885   0.7041305234645386   0.7012202358686404   0.1952797334681478   0.31502663691190286   0.8693346894522327   0.26770095227109536   0.44708183770837556   0.2529901428233342   0.543786247958635   0.3964491364695007   0.7427167034745258   0.7263101381353624   0.915405186148664   0.16136586525644378   0.005438452020016976   0.12274866392631935   0.5579484725556242   0.5434723932178696   0.8136485530718852   0.5782360305013308   0.12259070038941959   0.02564711590035852   0.7253091319667128   0.9574017997173423   0.41846017692488097   0.32442688003171816   0.5300293984985649   0.6423751628054395   0.5491254874726483   0.05672592776062283   0.08294756079018935   0.38938501998210523   0.005339239514013295   0.6602767912911222   0.34023085731566355   0.6630748818467429   0.08993405336534933   0.49891092603467835   0.3347924052956466   0.5403262179204236   0.5319855808097252   0.9554385328168088   0.5211438522237614   0.9620901874190928   0.4093948804203056   0.9297914169164503   0.7958347202570486   0.00468838770175051   0.9909347034954246   0.6053645368847321   0.26580532175848376   0.36231322489631107
0.44180921602277634   0.5486386091241093   0.1828577609682944   0.9729282049142058   0.436469976508763   0.8883618178329872   0.8426269036526308   0.30985332306746294   0.3465359231434137   0.3894508917983088   0.5078344983569844   0.7695271051470394   0.8145503423336885   0.4340123589815   0.986690646133223   0.8074369177279466   0.4051554619133829   0.5042209420650496   0.19085592587617434   0.8027485300261961   0.4142207584179583   0.8988564051803175   0.9250506041176906   0.44043530512988505   0.972411542395182   0.3502177960562083   0.7421928431493962   0.46750710021567926   0.535941565886419   0.46185597822322116   0.8995659394967653   0.15765377714821632   0.18940564274300523   0.07240508642491235   0.39173144113978103   0.3881266720011769   0.37485530040931675   0.6383927274434124   0.40504079500655804   0.5806897542732303   0.9696998384959338   0.13417178537836272   0.21418486913038373   0.7779412242470342   0.5554790800779755   0.23531538019804515   0.2891342650126931   0.33750591911714917   0.5830675376827935   0.8850975841418369   0.546941421863297   0.8699988189014699   0.04712597179637458   0.42324160591861576   0.6473754823665316   0.7123450417532536   0.8577203290533694   0.35083651949370337   0.2556440412267506   0.3242183697520767   0.4828650286440526   0.712443792050291   0.8506032462201926   0.7435286154788464
0.5131651901481188   0.5782720066719284   0.6364183770898089   0.9655873912318123   0.9576861100701434   0.34295662647388314   0.3472841120771157   0.628081472114663   0.3746185723873498   0.4578590423320463   0.8003426902138188   0.7580826532131931   0.32749260059097524   0.03461743641343054   0.15296720784728712   0.045737611459939514   0.46977227153760587   0.6837809169197272   0.8973231666205365   0.7215192417078629   0.9869072428935532   0.9713371248694361   0.04671992040034395   0.9779906262290164   0.47374205274543446   0.39306511819750783   0.41030154331053514   0.012403234997204199   0.5160559426752911   0.05010849172362471   0.06301743123341944   0.38432176288254116   0.14143737028794132   0.5922494493915784   0.2626747410196007   0.626239109669348   0.8139447696969662   0.5576320129781479   0.10970753317231358   0.5805014982094086   0.34417249815936024   0.8738510960584207   0.2123843665517771   0.8589822565015457   0.357265255265807   0.9025139711889846   0.1656644461514331   0.8809916302725294   0.8835232025203725   0.5094488529914767   0.755362902840898   0.868588395275325   0.36746725984508144   0.45934036126785205   0.6923454716074786   0.48426663239278395   0.22602988955714012   0.8670909118762736   0.42967073058787786   0.858027522723436   0.412085119860174   0.3094588988981257   0.3199631974155643   0.2775260245140274
0.06791262170081376   0.43560780283970496   0.10757883086378721   0.4185437680124817   0.7106473664350068   0.5330938316507204   0.9419143847123541   0.5375521377399524   0.8271241639146342   0.023644978659243667   0.1865514818714561   0.6689637424646273   0.4596569040695528   0.5643046173913916   0.49420601026397754   0.18469711007184333   0.23362701451241263   0.6972137055151181   0.06453527967609966   0.3266695873484074   0.8215418946522386   0.38775480661699235   0.7445720822605354   0.04914356283438001   0.7536292729514249   0.9521470037772873   0.6369932513967481   0.6305997948218983   0.042981906516418096   0.41905317212656695   0.6950788666843941   0.09304765708194593   0.2158577426017839   0.3954081934673233   0.508527384812938   0.42408391461731865   0.7562008385322311   0.8311035760759317   0.014321374548960462   0.2393868045454753   0.5225738240198184   0.1338898705608136   0.9497860948728608   0.9127172171970679   0.7010319293675799   0.7461350639438212   0.2052140126123254   0.8635736543626878   0.947402656416155   0.7939880601665339   0.5682207612155773   0.23297385954078959   0.9044207498997369   0.37493488803996694   0.8731418945311832   0.13992620245884366   0.688563007297953   0.9795266945726436   0.36461450971824516   0.715842287841525   0.9323621687657219   0.14842311849671203   0.35029313516928473   0.4764554832960497
0.40978834474590337   0.014533247935898408   0.4005070402964239   0.5637382660989818   0.7087564153783236   0.26839818399207716   0.19529302768409848   0.7001646117362939   0.7613537589621686   0.4744101238255432   0.6270722664685212   0.4671907521955043   0.8569330090624317   0.09947523578557628   0.7539303719373381   0.3272645497366607   0.1683700017644787   0.11994854121293262   0.3893158622190929   0.6114222618951357   0.23600783299875683   0.9715254227162206   0.03902272704980821   0.13496677859908598   0.8262194882528534   0.9569921747803222   0.6385156867533843   0.5712285125001042   0.1174630728745299   0.688593990788245   0.4432226590692858   0.8710639007638104   0.35610931391236134   0.21418386696270184   0.8161503926007646   0.403873148568306   0.49917630484992964   0.11470863117712556   0.062220020663426474   0.07660859883164532   0.33080630308545095   0.994760089964193   0.6729041584443336   0.4651863369365096   0.09479847008669408   0.023234667247972334   0.6338814313945254   0.33021955833742367   0.26857898183384066   0.06624249246765014   0.995365744641141   0.7589910458373195   0.15111590895931074   0.37764850167940506   0.5521430855718552   0.8879271450735091   0.7950065950469494   0.16346463471670325   0.7359926929710906   0.48405399650520314   0.2958302901970198   0.0487560035395777   0.6737726723076641   0.4074453976735578
0.9650239871115689   0.05399591357538477   0.0008685138633306242   0.9422590607370481   0.8702255170248748   0.030761246327412433   0.3669870824688053   0.6120395023996245   0.6016465351910342   0.9645187538597623   0.37162133782766427   0.8530484565623051   0.4505306262317234   0.5868702521803573   0.8194782522558091   0.965121311488796   0.655524031184774   0.42340561746365396   0.08348555928471837   0.48106731498359284   0.35969374098775425   0.37464961392407625   0.4097128869770542   0.07362191731003505   0.39466975387618536   0.3206537003486915   0.40884437311372357   0.13136285657298688   0.5244442368513106   0.28989245402127906   0.04185729064491829   0.5193233541733624   0.9227977016602764   0.3253737001615168   0.670235952817254   0.6662748976110573   0.472267075428553   0.7385034479811595   0.850757700561445   0.7011535861222613   0.816743044243779   0.3150978305175056   0.7672721412767266   0.2200862711386685   0.4570493032560248   0.9404482165934294   0.35755925429967245   0.14646435382863343   0.06237954937983943   0.6197945162447378   0.9487148811859488   0.015101497255646548   0.5379353125285289   0.3299020622234588   0.9068575905410305   0.4957781430822842   0.6151376108682524   0.004528362061942015   0.23662163772377653   0.8295032454712269   0.14287053543969938   0.2660249140807825   0.3858639371623315   0.12834965934896553
0.3261274911959203   0.9509270835632769   0.6185917958856049   0.9082633882102971   0.8690781879398956   0.010478866969847544   0.2610325415859325   0.7617990343816636   0.8066986385600561   0.3906843507251097   0.3123176603999836   0.746697537126017   0.2687633260315273   0.060782288501650926   0.405460069858953   0.25091939404373287   0.6536257151632748   0.05625392643970891   0.1688384321351765   0.42141614857250603   0.5107551797235755   0.7902290123589264   0.782974494972845   0.2930664892235405   0.18462768852765515   0.8393019287956496   0.16438269908724004   0.38480310101324344   0.3155495005877596   0.828823061825802   0.9033501575013075   0.6230040666315798   0.5088508620277035   0.4381387111006923   0.591032497101324   0.8763065295055628   0.24008753599617622   0.3773564225990414   0.18557242724237097   0.6253871354618299   0.5864618208329013   0.3211024961593325   0.016733995107194474   0.20397098688932389   0.07570664110932582   0.530873483800406   0.2337595001343495   0.9109044976657834   0.8910789525816707   0.6915715550047564   0.06937680104710947   0.52610139665254   0.575529451993911   0.8627484931789544   0.16602664354580188   0.9030973300209602   0.06667858996620758   0.4246097820782621   0.5749941464444779   0.0267908005153973   0.8265910539700314   0.047253359479220734   0.38942171920210694   0.4014036650535674
0.24012923313713005   0.7261508633198882   0.37268772409491246   0.1974326781642435   0.16442259202780424   0.1952773795194822   0.13892822396056292   0.28652818049846007   0.27334363944613355   0.5037058245147258   0.06955142291345347   0.7604267838459201   0.6978141874522225   0.6409573313357713   0.9035247793676516   0.8573294538249601   0.6311355974860149   0.21634754925750918   0.3285306329231737   0.8305386533095628   0.8045445435159836   0.16909418977828844   0.9391089137210668   0.42913498825599533   0.5644153103788535   0.4429433264584002   0.5664211896261543   0.23170231009175185   0.39999271835104927   0.24766594693891797   0.42749296566559136   0.9451741295932917   0.1266490789049157   0.7439601224241922   0.3579415427521379   0.18474734574737162   0.4288348914526932   0.10300279108842092   0.45441676338448633   0.32741789192241155   0.7976992939666783   0.8866552418309117   0.1258861304613126   0.49687923861284883   0.9931547504506947   0.7175610520526233   0.18677721674024583   0.06774425035685346   0.4287394400718412   0.2746177255942231   0.6203560271140915   0.8360419402651016   0.028746721720791974   0.0269517786553051   0.19286306144850016   0.8908678106718099   0.9020976428158762   0.2829916562311129   0.8349215186963622   0.7061204649244383   0.4732627513631831   0.17998886514269197   0.38050475531187594   0.3787025730020267
0.6755634573965048   0.29333362331178026   0.25461862485056336   0.8818233343891778   0.6824087069458101   0.5757725712591569   0.0678414081103175   0.8140790840323244   0.25366926687396885   0.3011548456649339   0.447485380996226   0.9780371437672228   0.22492254515317686   0.27420306700962876   0.2546223195477258   0.08716933309541294   0.3228249023373006   0.9912114107785159   0.4197008008513635   0.3810488681709747   0.8495621509741175   0.811222545635824   0.039196045539487585   0.0023462951689480318   0.1739986935776127   0.5178889223240437   0.7845774206889242   0.12052296077977018   0.4915899866318026   0.9421163510648868   0.7167360125786068   0.3064438767474458   0.23792071975783377   0.6409615053999529   0.2692506315823808   0.328406732980223   0.0129981746046569   0.36675843839032407   0.01462831203465496   0.24123739988481005   0.6901732722673564   0.3755470276118082   0.5949275111832915   0.8601885317138354   0.8406111212932388   0.5643244819759843   0.5557314656438038   0.8578422365448873   0.6666124277156261   0.04643555965194056   0.7711540449548796   0.7373192757651171   0.1750224410838235   0.1043192085870538   0.05441803237627286   0.43087539901767136   0.9371017213259897   0.46335770318710096   0.7851674007938921   0.10246866603744836   0.9241035467213328   0.09659926479677684   0.7705390887592372   0.8612312661526383
0.23393027445397652   0.7210522371849687   0.17561157757594573   0.001042734438802988   0.39331915316073773   0.15672775520898438   0.6198801119321419   0.14320049789391567   0.7267067254451116   0.11029219555704382   0.8487260669772623   0.40588122212879857   0.5516842843612881   0.005972986969990006   0.7943080346009894   0.9750058231111272   0.6145825630352983   0.542615283782889   0.009140633807097332   0.8725371570736788   0.6904790163139656   0.4460160189861122   0.2386015450478602   0.011305890921040512   0.45654874185998906   0.7249637818011436   0.06298996747191449   0.010263156482237523   0.06322958869925134   0.5682360265921592   0.4431098555397726   0.8670626585883219   0.3365228632541397   0.4579438310351154   0.5943837885625103   0.4611814364595233   0.7848385788928516   0.4519708440651254   0.8000757539615209   0.4861756133483961   0.17025601585755323   0.9093555602822363   0.7909351201544236   0.6136384562747172   0.47977699954358766   0.4633395412961241   0.5523335751065633   0.6023325653536767   0.023228257683598628   0.7383757594949805   0.48934360763464885   0.5920694088714392   0.9599986689843473   0.1701397329028213   0.04623375209487627   0.7250067502831173   0.6234758057302076   0.7121959018677059   0.45184996353236595   0.2638253138235941   0.838637226837356   0.26022505780258054   0.6517742095708451   0.777649700475198
0.6683812109798026   0.35086949752034424   0.8608390894164215   0.16401124420048077   0.188604211436215   0.8875299562242202   0.3085055143098581   0.561678678846804   0.16537595375261638   0.14915419672923963   0.8191619066752093   0.9696092699753648   0.20537728476826908   0.9790144638264183   0.772928154580333   0.24460251969224744   0.5819014790380616   0.2668185619587124   0.32107819104796703   0.9807772058686534   0.7432642522007056   0.00659350415613189   0.669303981477122   0.20312750539345534   0.07488304122090292   0.6557240066357877   0.8084648920607005   0.03911626119297459   0.886278829784688   0.7681940504115675   0.49995937775084237   0.47743758234617056   0.7209028760320716   0.619039853682328   0.6807974710756332   0.5078283123708057   0.5155255912638025   0.6400253898559096   0.9078693164953001   0.26322579267855833   0.9336241122257409   0.37320682789719717   0.586791125447333   0.282448586809905   0.19035986002503533   0.36661332374106526   0.917487143970211   0.07932108141644961   0.1154768188041324   0.7108893171052776   0.10902225190951059   0.04020482022347503   0.22919798901944446   0.9426952666937101   0.6090628741586682   0.5627672378773044   0.508295112987373   0.3236554130113821   0.9282654030830351   0.05493892550649871   0.9927695217235705   0.6836300231554726   0.020396086587735007   0.7917131328279404
0.05914540949782954   0.3104231952582754   0.4336049611404019   0.5092645460180354   0.8687855494727942   0.9438098715172101   0.5161178171701909   0.42994346460158583   0.7533087306686618   0.23292055441193252   0.40709556526068025   0.3897386443781108   0.5241107416492173   0.2902252877182224   0.798032691102012   0.8269714065008064   0.015815628661844407   0.9665698747068403   0.869767288018977   0.7720324809943077   0.023046106938273938   0.28293985155136775   0.8493712014312419   0.9803193481663672   0.9639006974404444   0.9725166562930924   0.41576624029084   0.4710548021483318   0.0951151479676502   0.02870678477588224   0.8996484231206491   0.041111337546745966   0.34180641729898836   0.7957862303639497   0.4925528578599689   0.6513726931686352   0.8176956756497711   0.5055609426457273   0.6945201667579568   0.8244012866678289   0.8018800469879266   0.538991067938887   0.8247528787389798   0.05236880567352127   0.7788339400496527   0.25605121638751926   0.975381677307738   0.07204945750715407   0.8149332426092083   0.2835345600944269   0.559615437016898   0.6009946553588222   0.7198180946415581   0.25482777531854467   0.6599670138962489   0.5598833178120763   0.37801167734256974   0.4590415449545949   0.16741415603628   0.9085106246434411   0.5603160016927987   0.9534806023088677   0.47289398927832316   0.08410933797561225
0.758435954704872   0.41448953436998065   0.6481411105393433   0.03174053230209098   0.9796020146552193   0.15843831798246139   0.6727594332316054   0.9596910747949369   0.16466877204601107   0.8749037578880345   0.11314399621470732   0.35869641943611463   0.444850677404453   0.6200759825694898   0.4531769823184585   0.7988131016240383   0.06683900006188326   0.1610344376148949   0.2857628262821785   0.8903024769805972   0.5065229983690845   0.20755383530602728   0.8128688370038553   0.8061931390049849   0.7480870436642125   0.7930643009360466   0.164727726464512   0.774452606702894   0.7684850290089932   0.6346259829535853   0.4919682932329067   0.8147615319079571   0.603816256962982   0.7597222250655508   0.37882429701819936   0.4560651124718424   0.15896557955852908   0.13964624249606095   0.9256473146997409   0.657252010847804   0.09212657949664582   0.9786118048811661   0.6398844884175624   0.7669495338672069   0.5856035811275613   0.7710579695751387   0.8270156514137071   0.960756394862222   0.8375165374633488   0.9779936686390921   0.6622879249491951   0.18630378815932797   0.06903150845435559   0.3433676856855069   0.17031963171628842   0.37154225625137094   0.46521525149137355   0.5836454606199561   0.7914953346980891   0.9154771437795285   0.30624967193284447   0.4439992181238952   0.8658480199983482   0.25822513293172444
0.21412309243619865   0.46538741324272914   0.22596353158078566   0.49127559906451757   0.6285195113086374   0.6943294436675904   0.39894788016707855   0.5305192042022956   0.7910029738452886   0.7163357750284982   0.7366599552178834   0.3442154160429676   0.721971465390933   0.37296808934299136   0.566340323501595   0.9726731597915967   0.25675621389955955   0.7893226287230353   0.7748449888035059   0.05719601601206821   0.950506541966715   0.34532341059914   0.9089969688051578   0.7989708830803438   0.7363834495305165   0.8799359973564108   0.6830334372243722   0.30769528401582624   0.10786393822187904   0.18560655368882048   0.2840855570572936   0.7771760798135307   0.3168609643765904   0.4692707786603222   0.5474256018394102   0.43296066377056297   0.5948894989856574   0.09630268931733085   0.9810852783378152   0.46028750397896623   0.33813328508609775   0.3069800605942956   0.20624028953430928   0.40309148796689803   0.38762674311938267   0.9616566499951555   0.29724332072915144   0.6041206048865543   0.6512432935888662   0.08172065263874473   0.6142098835047793   0.29642532087072804   0.5433793553669872   0.8961140989499242   0.3301243264474857   0.5192492410571974   0.22651839099039683   0.42684332028960204   0.7826987246080754   0.08628857728663444   0.6316288920047396   0.3305406309722712   0.8016134462702602   0.6260010733076682
0.2934956069186418   0.02356057037797557   0.5953731567359509   0.22290958534077016   0.9058688637992591   0.06190392038281998   0.2981298360067995   0.6187889804542159   0.25462557021039284   0.9801832677440753   0.6839199525020202   0.32236365958348784   0.7112462148434057   0.084069168794151   0.3537956260545345   0.8031144185262904   0.4847278238530088   0.6572258485045489   0.571096901446459   0.716825841239656   0.8530989318482692   0.32668521753227775   0.7694834551761988   0.09082476793198777   0.5596033249296275   0.3031246471543022   0.1741102984402478   0.8679151825912176   0.6537344611303684   0.2412207267714822   0.8759804624334483   0.24912620213700173   0.39910889091997553   0.26103745902740694   0.19206050993142812   0.9267625425535139   0.6878626760765699   0.17696829023325597   0.8382648838768936   0.12364812402722347   0.20313485222356112   0.519742441728707   0.2671679824304346   0.4068222827875675   0.3500359203752919   0.19305722419642926   0.49768452725423584   0.31599751485557975   0.7904325954456645   0.889932577042127   0.323574228813988   0.4480823322643621   0.1366981343152961   0.6487118502706448   0.4475937663805397   0.19895613012736038   0.7375892433953206   0.3876743912432379   0.25553325644911157   0.2721935875738465   0.049726567318750664   0.21070610100998194   0.41726837257221794   0.148545463546623
0.8465917150951895   0.6909636592812749   0.15010039014178334   0.7417231807590555   0.49655579471989764   0.49790643508484567   0.6524158628875475   0.42572566590347577   0.7061231992742332   0.6079738580427186   0.3288416340735595   0.9776433336391136   0.5694250649589371   0.9592620077720737   0.8812478676930198   0.7786872035117532   0.8318358215636166   0.5715876165288358   0.6257146112439083   0.5064936159379068   0.7821092542448659   0.36088151551885395   0.20844623867169032   0.35794815239128375   0.9355175391496763   0.669917856237579   0.05834584852990698   0.6162249716322282   0.4389617444297787   0.17201142115273335   0.4059299856423595   0.19049930572875248   0.7328385451555455   0.5640375631100147   0.07708835156879996   0.21285597208963886   0.16341348019660842   0.604775555337941   0.19584048387578015   0.4341687685778856   0.3315776586329919   0.03318793880910512   0.5701258726318719   0.9276751526399788   0.549468404388126   0.6723064232902511   0.3616796339601816   0.569727000248695   0.6139508652384497   0.0023885670526721603   0.3033337854302746   0.9535020286164668   0.174989120808671   0.8303771458999388   0.8974037997879152   0.7630027228877143   0.4421505756531255   0.26633958278992403   0.8203154482191152   0.5501467507980755   0.27873709545651704   0.6615640274519831   0.624474964343335   0.11597798222018989
0.9471594368235252   0.628376088642878   0.05434909171146312   0.18830282958021108   0.39769103243539916   0.9560696653526267   0.6926694577512815   0.618575829331516   0.7837401671969495   0.9536810982999546   0.3893356723210069   0.6650738007150492   0.6087510463882785   0.1233039524000158   0.49193187253309173   0.9020710778273349   0.166600470735153   0.8569643696100917   0.6716164243139766   0.3519243270292594   0.8878633752786359   0.19540034215810867   0.047141459970641536   0.2359463448090695   0.9407039384551108   0.5670242535152307   0.9927923682591784   0.04764351522885842   0.5430129060197116   0.610954588162604   0.3001229105078969   0.4290676858973424   0.7592727388227621   0.6572734898626493   0.91078723818689   0.7639938851822933   0.15052169243448366   0.5339695374626335   0.4188553656537983   0.8619228073549584   0.9839212216993306   0.6770051678525418   0.7472389413398217   0.5099984803256989   0.09605784642069472   0.48160482569443314   0.7000974813691802   0.2740521355166295   0.15535390796558393   0.9145805721792024   0.7073051131100018   0.22640862028777106   0.6123410019458724   0.30362598401659846   0.40718220260210486   0.7973409343904286   0.8530682631231101   0.6463524941539491   0.49639496441521486   0.03334704920813541   0.7025465706886265   0.1123829566913156   0.0775395987614166   0.17142424185317706
0.7186253489892959   0.4353777888387738   0.3303006574215949   0.6614257615274781   0.6225675025686012   0.9537729631443407   0.6302031760524147   0.3873736260108486   0.4672135946030172   0.039192390965138275   0.922898062942413   0.16096500572307754   0.8548725926571449   0.7355664069485398   0.5157158603403081   0.3636240713326489   0.0018043295340346957   0.08921391279459068   0.01932089592509333   0.3302770221245135   0.2992577588454082   0.9768309561032751   0.9417812971636768   0.15885278027133645   0.5806324098561123   0.5414531672645013   0.6114806397420818   0.49742701874385836   0.9580649072875111   0.5876802041201606   0.9812774636896671   0.11005339273300978   0.49085131268449395   0.5484878131550223   0.05837940074725403   0.9490883870099323   0.6359787200273491   0.8129214062064825   0.5426635404069459   0.5854643156772833   0.6341743904933144   0.7237074934118918   0.5233426444818525   0.2551872935527698   0.3349166316479062   0.7468765373086167   0.5815613473181758   0.09633451328143335   0.7542842217917939   0.20542337004411546   0.970080707576094   0.598907494537575   0.7962193145042827   0.6177431659239548   0.9888032438864269   0.4888541018045652   0.30536800181978874   0.06925535276893256   0.9304238431391729   0.539765714794633   0.6693892817924397   0.25633394656245007   0.38776030273222706   0.9543013991173497
0.035214891299125285   0.5326264531505582   0.8644176582503745   0.6991141055645799   0.7002982596512191   0.7857499158419415   0.2828563109321987   0.6027795922831465   0.9460140378594252   0.580326545797826   0.31277560335610477   0.00387209774557152   0.14979472335514246   0.9625833798738712   0.32397235946967784   0.5150179959410064   0.8444267215353537   0.8933280271049386   0.39354851633050497   0.9752522811463734   0.17503743974291402   0.6369940805424885   0.005788213598277907   0.020950882029023742   0.13982254844378872   0.10436762739193031   0.14137055534790338   0.3218367764644439   0.43952428879256966   0.3186177115499888   0.8585142444157047   0.7190571841812974   0.4935102509331445   0.7382911657521628   0.5457386410595999   0.7151850864357259   0.343715527578002   0.7757077858782916   0.22176628158992207   0.20016709049471956   0.49928880604264836   0.882379758773353   0.8282177652594171   0.22491480934834618   0.32425136629973433   0.24538567823086438   0.8224295516611392   0.20396392731932245   0.18442881785594561   0.14101805083893407   0.6810589963132359   0.8821271508548786   0.7449045290633759   0.8224003392889453   0.8225447518975312   0.16306996667358112   0.25139427813023146   0.0841091735367825   0.2768061108379313   0.4478848802378552   0.9076787505522295   0.30840138765849096   0.055039829248009216   0.24771778974313566
0.4083899445095811   0.426021628885138   0.22682206398859212   0.022802980394789462   0.08413857820984677   0.18063595065427362   0.40439251232745294   0.818839053075467   0.8997097603539012   0.03961789981533958   0.7233335160142171   0.9367119022205885   0.15480523129052523   0.21721756052639432   0.900788764116686   0.7736419355470073   0.9034109531602937   0.13310838698961183   0.6239826532787547   0.32575705530915217   0.9957322026080643   0.8247069993311209   0.5689428240307455   0.07803926556601651   0.5873422580984832   0.3986853704459829   0.34212076004215336   0.05523628517122704   0.5032036798886365   0.21804941979170925   0.9377282477147004   0.23639723209576002   0.6034939195347353   0.17843151997636966   0.21439473170048332   0.29968532987517155   0.44868868824421004   0.9612139594499753   0.3136059675837974   0.5260433943281642   0.5452777350839163   0.8281055724603635   0.6896233143050428   0.20028633901901202   0.549545532475852   0.003398573129242641   0.12068049027429725   0.12224707345299553   0.9622032743773687   0.6047132026832598   0.7785597302321439   0.06701078828176849   0.45899959448873234   0.3866637828915505   0.8408314825174434   0.8306135561860084   0.8555056749539971   0.20823226291518082   0.6264367508169602   0.5309282263108369   0.40681698670978705   0.24701830346520548   0.31283078323316277   0.004884831982672729
0.8615392516258708   0.41891273100484194   0.6232074689281201   0.8045984929636607   0.3119937191500188   0.4155141578755993   0.5025269786538228   0.6823514195106651   0.34979044477265   0.8108009551923395   0.7239672484216789   0.6153406312288967   0.8907908502839177   0.42413717230078907   0.8831357659042355   0.7847270750428882   0.035285175329920586   0.21590490938560822   0.2566990150872753   0.25379884873205133   0.6284681886201335   0.9688866059204028   0.9438682318541125   0.24891401674937857   0.7669289369942628   0.5499738749155608   0.32066076292599244   0.44431552378571787   0.45493521784424407   0.13445971703996146   0.8181337842721697   0.7619641042750527   0.10514477307159405   0.32365876184762193   0.09416653585049072   0.14662347304615603   0.2143539227876764   0.8995215895468328   0.21103076994625528   0.36189639800326784   0.1790687474577558   0.6836166801612247   0.95433175485898   0.10809754927121651   0.5506005588376223   0.7147300742408219   0.010463523004867494   0.859183532521838   0.7836716218433595   0.16475619932526114   0.6898027600788751   0.41486800873612006   0.32873640399911536   0.03029648228529967   0.8716689758067054   0.6529039044610674   0.22359163092752132   0.7066377204376778   0.7775024399562147   0.5062804314149113   0.009237708139844949   0.8071161308908449   0.5664716700099595   0.1443840334116435
0.8301689606820891   0.12349945072962025   0.6121399151509794   0.036286484140426976   0.2795684018444669   0.40876937648879835   0.6016763921461119   0.17710295161858905   0.4958967800011075   0.2440131771635372   0.9118736320672369   0.762234942882469   0.1671603760019921   0.21371669487823752   0.04020465626053146   0.10933103842140166   0.9435687450744707   0.5070789744405598   0.2627022163043167   0.6030506070064904   0.9343310369346258   0.6999628435497148   0.6962305462943573   0.45866657359484686   0.10416207625253666   0.5764633928200946   0.08409063114337784   0.42238008945441985   0.8245936744080697   0.1676940163312963   0.4824142389972659   0.24527713783583083   0.32869689440696226   0.9236808391677591   0.570540606930029   0.4830421949533618   0.16153651840497016   0.7099641442895216   0.5303359506694976   0.3737111565319602   0.21796777333049938   0.20288516984896177   0.2676337343651808   0.7706605495254698   0.28363673639587356   0.5029223262992469   0.5714031880708235   0.311993975930623   0.1794746601433369   0.9264589334791523   0.48731255692744563   0.8896138864762031   0.35488098573526716   0.758764917147856   0.004898317930179765   0.6443367486403723   0.026184091328304893   0.8350840779800969   0.4343577110001508   0.16129455368701046   0.8646475729233347   0.12511993369057536   0.9040217603306533   0.7875833971550502
0.6466797995928354   0.9222347638416136   0.6363880259654725   0.01692284762958041   0.3630430631969618   0.4193124375423667   0.06498483789464898   0.7049288716989575   0.18356840305362485   0.49285350406321443   0.5776722809672034   0.8153149852227544   0.8286874173183577   0.7340885869153584   0.5727739630370235   0.17097823658238204   0.8025033259900528   0.8990045089352615   0.1384162520368728   0.009683682895371583   0.9378557530667181   0.7738845752446861   0.23439449170621954   0.22210028574032134   0.29117595347388275   0.8516498114030726   0.598006465740747   0.20517743811074093   0.9281328902769209   0.43233737386070586   0.5330216278460981   0.5002485664117835   0.7445644872232962   0.9394838697974914   0.9553493468788947   0.6849335811890291   0.9158770699049384   0.20539528288213302   0.3825753838418712   0.5139553446066472   0.11337374391488562   0.3063907739468715   0.24415913180499837   0.5042716617112756   0.17551799084816755   0.5325061987021853   0.009764640098778832   0.28217137597095426   0.8843420373742849   0.6808563872991127   0.4117581743580318   0.07699393786021333   0.9562091470973638   0.24851901343840685   0.8787365465119337   0.5767453714484299   0.21164465987406772   0.3090351436409154   0.923387199633039   0.8918117902594006   0.2957675899691293   0.10363986075878236   0.5408118157911678   0.37785644565275345
0.18239384605424366   0.7972490868119109   0.29665268398616945   0.8735847839414779   0.006875855206076121   0.26474288810972557   0.28688804388739064   0.5914134079705237   0.1225338178317913   0.5838865008106129   0.8751298695293589   0.5144194701103103   0.16632467073442747   0.335367487372206   0.9963933230174251   0.9376740986618805   0.9546800108603597   0.026332343731290633   0.07300612338438615   0.04586230840247983   0.6589124208912305   0.9226924829725083   0.5321943075932184   0.6680058627497264   0.4765185748369868   0.12544339616059738   0.2355416236070489   0.7944210788082484   0.46964271963091064   0.8607005080508718   0.9486535797196582   0.20300767083772484   0.34710890179911935   0.27681400724025895   0.07352371019029942   0.6885882007274146   0.18078423106469188   0.941446519868053   0.07713038717287428   0.7509141020655341   0.22610422020433216   0.9151141761367623   0.004124263788488121   0.7050517936630543   0.5671917993131017   0.992421693164254   0.4719299561952698   0.037045930913327856   0.09067322447611495   0.8669782970036567   0.2363883325882209   0.2426248521050794   0.6210305048452043   0.0062777889527848366   0.28773475286856265   0.039617181267354556   0.273921603046085   0.7294637817125259   0.2142110426782632   0.35102898053994   0.09313737198139307   0.788017261844473   0.13708065550538892   0.600114878474406
0.867033151777061   0.8729030857077106   0.1329563917169008   0.8950630848113518   0.2998413524639592   0.8804813925434566   0.661026435521631   0.8580171538980239   0.2091681279878443   0.01350309553979991   0.42463810293341014   0.6153923017929445   0.58813762314264   0.007225306587015073   0.1369033500648475   0.57577512052559   0.314216020096555   0.2777615248744892   0.9226923073865843   0.22474613998564993   0.22107864811516195   0.4897442630300163   0.7856116518811954   0.6246312615112439   0.354045496338101   0.6168411773223057   0.6526552601642945   0.7295681766998922   0.05420414387414179   0.7363597847788491   0.9916288246426636   0.8715510228018682   0.8450360158862975   0.7228566892390492   0.5669907217092534   0.25615872100892373   0.2568983927436575   0.7156313826520341   0.4300873716444059   0.6803836004833338   0.9426823726471025   0.43786985777754495   0.5073950642578217   0.4556374604976839   0.7216037245319405   0.9481255947475287   0.7217834123766262   0.8310061989864399   0.36755822819383954   0.33128441742522297   0.06912815221233166   0.10143802228654776   0.31335408431969775   0.5949246326463739   0.07749932756966812   0.2298869994846795   0.46831806843340024   0.8720679434073246   0.5105086058604147   0.9737282784757557   0.21141967568974274   0.15643656075529055   0.08042123421600882   0.2933446779924219
0.2687373030426402   0.7185667029777456   0.5730261699581872   0.8377072174947381   0.5471335785106997   0.7704411082302169   0.851242757581561   0.006701018508298127   0.17957535031686012   0.439156690804994   0.7821146053692293   0.9052629962217503   0.8662212659971623   0.8442320581586201   0.7046152777995612   0.6753759967370709   0.39790319756376213   0.9721641147512955   0.19410667193914646   0.7016477182613151   0.18648352187401937   0.8157275539960049   0.11368543772313766   0.40830304026889325   0.9177462188313792   0.09716085101825929   0.5406592677649504   0.5705958227741552   0.3706126403206795   0.32671974278804233   0.6894165101833895   0.563894804265857   0.19103729000381936   0.8875630519830483   0.9073019048141602   0.6586318080441067   0.324816024006657   0.04333099382442819   0.202686627014599   0.9832558113070358   0.9269128264428949   0.07116687907313272   0.008579955075452521   0.2816080930457206   0.7404293045688756   0.2554393250771278   0.8948945173523148   0.8733050527768274   0.8226830857374964   0.15827847405886852   0.3542352495873644   0.30270923000267225   0.45207044541681685   0.8315587312708262   0.664818739403975   0.7388144257368152   0.2610331554129975   0.9439956792877778   0.7575168345898148   0.08018261769270854   0.9362171314063404   0.9006646854633497   0.5548302075752158   0.09692680638567278
0.009304304963445585   0.829497806390217   0.5462502524997632   0.8153187133399521   0.2688750003945701   0.5740584813130891   0.6513557351474484   0.9420136605631247   0.4461919146570737   0.41578000725422065   0.29712048556008397   0.6393044305604525   0.9941214692402568   0.5842212759833945   0.632301746156109   0.9004900048236373   0.7330883138272594   0.6402255966956165   0.8747849115662942   0.8203073871309288   0.7968711824209188   0.7395609112322669   0.3199547039910785   0.723380580745256   0.7875668774574732   0.9100631048420499   0.7737044514913152   0.9080618674053038   0.5186918770629032   0.33600462352896077   0.12234871634386682   0.9660482068421791   0.0724999624058295   0.9202246162747402   0.8252282307837828   0.3267437762817266   0.07837849316557266   0.3360033402913457   0.1929264846276738   0.4262537714580893   0.34529017933831335   0.6957777435957292   0.3181415730613795   0.6059463843271605   0.5484189969173945   0.9562168323634623   0.9981868690703011   0.8825658035819045   0.7608521194599213   0.0461537275214124   0.22448241757898585   0.9745039361766007   0.24216024239701806   0.7101491039924517   0.10213370123511903   0.008455729334421649   0.16966027999118857   0.7899244877177115   0.2769054704513362   0.681711953052695   0.09128178682561591   0.4539211474263658   0.08397898582366238   0.2554581815946058
0.7459916074873025   0.7581434038306367   0.7658374127622828   0.6495117972674452   0.19757261056990807   0.8019265714671744   0.7676505436919817   0.7669459936855407   0.43672049110998684   0.7557728439457619   0.5431681261129959   0.7924420575089399   0.19456024871296876   0.04562373995331033   0.44103442487787686   0.7839863281745183   0.02489996872178018   0.2556992522355988   0.16412895442654069   0.10227437512182326   0.9336181818961643   0.801778104809233   0.0801499686028783   0.8468161935272175   0.18762657440886168   0.04363470097859633   0.3143125558405955   0.1973043962597722   0.9900539638389536   0.24170812951142195   0.5466620121486138   0.43035840257423147   0.5533334727289668   0.48593528556565996   0.003493886035617822   0.6379163450652915   0.35877322401599804   0.44031154561234964   0.5624594611577409   0.8539300168907732   0.3338732552942179   0.18461229337675084   0.39833050673120024   0.75165564176895   0.4002550733980536   0.38283418856751783   0.318180538128322   0.9048394482417325   0.21262849898919192   0.3391994875889215   0.003867982287726466   0.7075350519819603   0.22257453515023828   0.09749135807749956   0.45720597013911274   0.2771766494077288   0.6692410624212715   0.6115560725118396   0.4537120841034949   0.6392603043424373   0.3104678384052734   0.17124452689948994   0.8912526229457539   0.7853302874516641
0.9765945831110555   0.9866322335227391   0.49292211621455373   0.03367464568271417   0.5763395097130019   0.6037980449552213   0.17474157808623175   0.1288351974409817   0.36371101072380996   0.2645985573662997   0.17087359579850528   0.42130014545902145   0.1411364755735717   0.1671071992888002   0.7136676256593926   0.14412349605129265   0.4718954131523002   0.5555511267769606   0.2599555415558976   0.5048631917088554   0.16142757474702682   0.3843065998774707   0.36870291861014365   0.7195329042571913   0.18483299163597128   0.3976743663547316   0.87578080239559   0.6858582585744771   0.6084934819229694   0.7938763213995103   0.7010392243093582   0.5570230611334954   0.2447824711991594   0.5292777640332106   0.5301656285108529   0.13572291567447395   0.10364599562558773   0.36217056474441034   0.8164980028514603   0.9915994196231813   0.6317505824732875   0.8066194379674497   0.5565424612955627   0.4867362279143259   0.4703230077262607   0.4223128380899791   0.18783954268541905   0.7672033236571346   0.2854900160902894   0.024638471735247535   0.3120587402898291   0.08134506508265754   0.67699653416732   0.23076215033573724   0.6110195159804709   0.5243220039491622   0.4322140629681606   0.7014843863025267   0.080853887469618   0.3885990882746882   0.3285680673425729   0.33931382155811635   0.2643558846181576   0.3969996686515069
0.6968174848692854   0.5326943835906666   0.7078134233225949   0.9102634407371809   0.22649447714302468   0.11038154550068749   0.5199738806371759   0.14306011708004632   0.9410044610527353   0.08574307376543995   0.20791514034734673   0.06171505199738876   0.26400792688541524   0.8549809234297027   0.5968956243668758   0.5373930480482266   0.8317938639172546   0.153496537127176   0.5160417368972579   0.1487939597735384   0.5032257965746818   0.8141827155690596   0.2516858522791002   0.7517942911220316   0.8064083117053964   0.2814883319783931   0.5438724289565053   0.8415308503848505   0.5799138345623718   0.1711067864777056   0.023898548319329464   0.6984707333048042   0.6389093735096365   0.08536371271226567   0.8159834079719828   0.6367556813074156   0.3749014466242212   0.23038278928256298   0.21908778360510692   0.0993626332591889   0.5431075827069666   0.07688625215538696   0.7030460467078491   0.9505686734856504   0.03988178613228481   0.2627035365863273   0.4513601944287489   0.19877438236361897   0.2334734744268884   0.9812152046079342   0.9074877654722436   0.3572435319787684   0.6535596398645167   0.8101084181302285   0.8835892171529142   0.6587727986739641   0.014650266354880204   0.7247447054179629   0.0676058091809314   0.022017117366548624   0.639748819730659   0.4943619161353999   0.8485180255758245   0.9226544841073597
0.0966412370236924   0.41747566398001296   0.1454719788679754   0.9720858106217093   0.05675945089140759   0.15477212739368568   0.6941117844392265   0.7733114282580903   0.8232859764645192   0.17355692278575152   0.7866240189669829   0.4160678962793219   0.1697263366000025   0.363448504655523   0.9030348018140687   0.7572950976053577   0.1550760702451223   0.6387037992375602   0.8354289926331373   0.7352779802388092   0.5153272505144634   0.1443418831021602   0.9869109670573128   0.8126234961314495   0.41868601349077095   0.7268662191221472   0.8414389881893375   0.8405376855097402   0.36192656259936334   0.5720940917284616   0.14732720375011102   0.06722625725164989   0.5386405861348441   0.3985371689427101   0.36070318478312813   0.651158360972328   0.36891424953484164   0.035088664287187064   0.45766838296905943   0.8938632633669702   0.21383817928971935   0.39638486504962694   0.6222393903359221   0.15858528312816106   0.698510928775256   0.25204298194746677   0.6353284232786092   0.34596178699671165   0.2798249152844851   0.5251767628253194   0.7938894350892717   0.5054241014869715   0.9178983526851218   0.953082671096858   0.6465622313391607   0.43819784423532154   0.3792577665502776   0.5545455021541479   0.28585904655603256   0.7870394832629936   0.010343517015435962   0.5194568378669608   0.8281906635869731   0.8931762198960234
0.7965053377257166   0.12307197281733386   0.2059512732510511   0.7345909367678622   0.09799440895046056   0.8710289908698671   0.5706228499724418   0.38862914977115065   0.8181694936659755   0.3458522280445476   0.7767334148831702   0.8832050482841792   0.9002711409808537   0.3927695569476897   0.13017118354400942   0.44500720404885763   0.521013374430576   0.8382240547935418   0.8443121369879768   0.6579677207858641   0.5106698574151401   0.318767216926581   0.01612147340100369   0.7647915008898407   0.7141645196894235   0.19569524410924719   0.8101702001499526   0.03020056412197839   0.6161701107389629   0.3246662532393801   0.23954735017751075   0.6415714143508278   0.7980006170729874   0.9788140251948324   0.4628139352943406   0.7583663660666485   0.8977294760921338   0.5860444682471427   0.3326427517503312   0.3133591620177909   0.3767161016615577   0.747820413453601   0.48833061476235434   0.6553914412319268   0.8660462442464176   0.4290531965270199   0.4722091413613506   0.8905999403420861   0.15188172455699414   0.23335795241777274   0.6620389412113981   0.8603993762201078   0.5357116138180312   0.9086916991783927   0.4224915910338873   0.21882796186928002   0.7377109967450437   0.9298776739835602   0.9596776557395467   0.4604615958026315   0.83998152065291   0.34383320573641746   0.6270349039892155   0.1471024337848406
0.4632654189913522   0.5960127922828166   0.13870428922686118   0.4917109925529138   0.5972191747449346   0.1669595957557966   0.6664951478655106   0.6011110522108276   0.44533745018794046   0.9336016433380239   0.004456206654112501   0.7407116759907199   0.9096258363699092   0.024909944159631225   0.5819646156202252   0.5218837141214399   0.1719148396248655   0.09503227017607102   0.6222869598806785   0.06142211831880832   0.33193331897195555   0.7511990644396536   0.995252055891463   0.9143196845339677   0.8686678999806033   0.15518627215683706   0.8565477666646019   0.42260869198105394   0.2714487252356687   0.9882266764010404   0.1900526187990913   0.8214976397702263   0.8261112750477283   0.05462503306301657   0.1855964121449788   0.08078596377950642   0.916485438677819   0.029715088903385343   0.6036317965247536   0.5589022496580666   0.7445705990529535   0.9346828187273143   0.9813448366440751   0.4974801313392583   0.412637280080998   0.18348375428766076   0.9860927807526121   0.5831604468052906   0.5439693801003946   0.028297482130823684   0.12954501408801022   0.16055175482423664   0.27252065486472593   0.040070805729783235   0.9394923952889189   0.33905411505401034   0.4464093798169977   0.9854457726667667   0.7538959831439401   0.2582681512745039   0.5299239411391787   0.9557306837633813   0.1502641866191865   0.6993659016164373
0.7853533420862252   0.02104786503606701   0.16891934997511143   0.20188577027717908   0.3727160620052272   0.8375641107484063   0.18282656922249937   0.6187253234718885   0.8287466819048326   0.8092666286175826   0.053281555134489164   0.45817356864765185   0.5562260270401066   0.7691958228877993   0.11378915984557025   0.1191194535936415   0.10981664722310891   0.7837500502210327   0.3598931767016302   0.8608513023191375   0.5798927060839302   0.8280193664576513   0.20962899008244365   0.16148540070270023   0.794539363997705   0.8069715014215844   0.040709640107332225   0.9595996304255211   0.4218233019924778   0.969407390673178   0.8578830708848328   0.34087430695363263   0.5930766200876452   0.1601407620555955   0.8046015157503437   0.8827007383059808   0.03685059304753859   0.39094493916779616   0.6908123559047734   0.7635812847123393   0.9270339458244297   0.6071948889467634   0.3309191792031433   0.9027299823932017   0.3471412397404995   0.7791755224891121   0.12129018912069962   0.7412445816905014   0.5526018757427944   0.9722040210675278   0.08058054901336739   0.7816449512649803   0.13077857375031665   0.0027966303943497447   0.22269747812853455   0.4407706443113477   0.5377019536626715   0.8426558683387543   0.41809596237819086   0.5580699060053669   0.5008513606151329   0.4517109291709581   0.7272836064734174   0.7944886212930277
0.5738174147907031   0.8445160402241947   0.39636442727027416   0.8917586388998259   0.2266761750502037   0.06534051773508251   0.27507423814957455   0.15051405720932443   0.6740742993074093   0.09313649666755469   0.19449368913620713   0.3688691059443441   0.5432957255570926   0.09033986627320495   0.9717962110076726   0.9280984616329964   0.005593771894421163   0.2476839979344507   0.5537002486294818   0.3700285556276295   0.5047424112792883   0.7959730687634926   0.8264166421560644   0.5755399343346018   0.9309249964885852   0.9514570285392979   0.43005221488579015   0.683781295434776   0.7042488214383814   0.8861165108042154   0.15497797673621563   0.5332672382254515   0.030174522130972128   0.7929800141366607   0.9604842876000085   0.16439813228110742   0.4868787965738795   0.7026401478634557   0.9886880765923359   0.23629967064811103   0.48128502467945833   0.45495614992900507   0.4349878279628542   0.8662711150204816   0.97654261340017   0.6589830811655125   0.6085711858067898   0.2907311806858797   0.045617616911584925   0.7075260526262146   0.1785189709209997   0.6069498852511038   0.34136879547320353   0.8214095418219992   0.023540994184784076   0.07368264702565229   0.3111942733422314   0.02842952768533842   0.0630567065847756   0.9092845147445449   0.8243154767683519   0.3257893798218826   0.07436862999243969   0.6729848440964339
0.34303045208889354   0.8708332298928776   0.6393808020295856   0.8067137290759523   0.3664878386887235   0.21185014872736502   0.03080961622279568   0.5159825483900726   0.3208702217771386   0.5043240961011505   0.852290645301796   0.9090326631389688   0.979501426303935   0.6829145542791513   0.8287496511170119   0.8353500161133165   0.6683071529617036   0.6544850265938128   0.7656929445322364   0.9260655013687716   0.8439916761933518   0.3286956467719302   0.6913243145397966   0.25308065727233775   0.5009612241044582   0.45786241687905266   0.051943512510211086   0.44636692819638546   0.13447338541573475   0.24601226815168767   0.02113389628741541   0.9303843798063128   0.8136031636385962   0.7416881720505373   0.16884325098561942   0.021351716667344058   0.8341017373346612   0.05877361777138597   0.34009359986860754   0.18600170055402754   0.16579458437295752   0.4042885911775731   0.5744006553363712   0.2599361991852559   0.3218029081796057   0.0755929444056429   0.8830763407965746   0.006855541912918152   0.8208416840751475   0.6177305275265902   0.8311328282863635   0.5604886137165327   0.6863682986594127   0.37171825937490255   0.8099989319989481   0.6301042339102199   0.8727651350208165   0.6300300873243654   0.6411556810133286   0.6087525172428758   0.0386633976861554   0.5712564695529794   0.30106208114472116   0.42275081668884823
0.8728688133131979   0.16696787837540625   0.7266614258083499   0.1628146175035923   0.5510659051335921   0.09137493396976333   0.8435850850117753   0.15595907559067415   0.7302242210584446   0.47364440644317307   0.012452256725411823   0.5954704618741414   0.043855922399031896   0.10192614706827052   0.20245332472646374   0.9653662279639216   0.17109078737821534   0.4718960597439052   0.5612976437131351   0.35661371072104586   0.13242738969205994   0.9006395901909259   0.2602355625684139   0.9338628940321977   0.25955857637886204   0.7336717118155196   0.533574136760064   0.7710482765286053   0.7084926712452699   0.6422967778457562   0.6899890517482887   0.6150892009379312   0.9782684501868253   0.16865237140258318   0.6775367950228769   0.019618739063789737   0.9344125277877934   0.06672622433431265   0.4750834702964131   0.05425251109986811   0.763321740409578   0.5948301645904075   0.9137858265832781   0.6976388003788222   0.6308943507175181   0.6941905743994816   0.6535502640148642   0.7637759063466246   0.37133577433865605   0.960518862583962   0.11997612725480013   0.9927276298180193   0.6628431030933861   0.3182220847382058   0.42998707550651144   0.3776384288800881   0.6845746529065608   0.14956971333562258   0.7524502804836346   0.35801968981629834   0.7501621251187675   0.08284348900130994   0.2773668101872215   0.3037671787164302
0.9868403847091894   0.4880133244109025   0.3635809836039434   0.606128378337608   0.35594603399167135   0.7938227500114209   0.7100307195890793   0.8423524719909834   0.9846102596530153   0.8333038874274589   0.5900545923342791   0.8496248421729641   0.3217671565596292   0.5150818026892531   0.16006751682776768   0.471986413292876   0.6371925036530683   0.3655120893536305   0.4076172363441331   0.11396672347657766   0.8870303785343009   0.28266860035232055   0.1302504261569116   0.8101995447601474   0.9001899938251114   0.794655275941418   0.7666694425529682   0.20407116642253945   0.5442439598334401   0.0008325259299971986   0.05663872296388891   0.3617186944315561   0.5596337001804248   0.16752863850253838   0.46658413062960974   0.5120938522585919   0.23786654362079562   0.6524468358132853   0.3065166138018421   0.04010743896571597   0.6006740399677273   0.28693474645965483   0.898899377457709   0.9261407154891383   0.7136436614334264   0.00426614610733431   0.7686489513007974   0.11594117072899089   0.813453667608315   0.20961087016591626   0.001979508747829202   0.9118700043064515   0.26920970777487485   0.20877834423591907   0.9453407857839403   0.5501513098748954   0.70957600759445   0.04124970573338068   0.4787566551543305   0.03805745761630342   0.4717094639736544   0.3888028699200954   0.17224004135248844   0.9979500186505874
0.8710354240059272   0.10186812346044052   0.27334066389477946   0.07180930316144914   0.1573917625725007   0.09760197735310622   0.504691712593982   0.9558681324324583   0.34393809496418576   0.88799110718719   0.5027122038461529   0.043998128126006786   0.07472838718931091   0.6792127629512709   0.5573714180622126   0.4938468182511114   0.36515237959486085   0.6379630572178903   0.07861476290788204   0.45578936063480796   0.8934429156212065   0.24916018729779485   0.9063747215553936   0.45783934198422055   0.022407491615279364   0.14729206383735433   0.6330340576606142   0.38603003882277137   0.8650157290427787   0.04969008648424811   0.12834234506663209   0.43016190639031315   0.5210776340785929   0.16169897929705815   0.6256301412204792   0.38616377826430637   0.446349246889282   0.48248621634578726   0.06825872315826664   0.8923169600131949   0.08119686729442113   0.844523159127897   0.9896439602503846   0.436527599378387   0.18775395167321465   0.5953629718301022   0.083269238694991   0.9786882573941664   0.1653464600579353   0.44807090799274785   0.4502351810343769   0.5926582185713951   0.3003307310151566   0.3983808215084998   0.3218928359677448   0.16249631218108193   0.7792530969365637   0.23668184221144162   0.6962626947472655   0.7763325339167756   0.3329038500472817   0.7541956258656544   0.6280039715889989   0.8840155739035807
0.2517069827528606   0.9096724667377574   0.6383600113386143   0.4474879745251936   0.06395303107964591   0.31430949490765514   0.5550907726436234   0.46879971713102714   0.8986065710217106   0.8662385869149073   0.10485559160924648   0.8761414985596321   0.598275840006554   0.4678577654064075   0.7829627556415018   0.7136451863785501   0.8190227430699902   0.23117592319496585   0.08670006089423613   0.9373126524617745   0.48611889302270855   0.4769802973293115   0.4586960893052372   0.05329707855819396   0.23441191026984798   0.5673078305915542   0.8203360779666228   0.6058091040330004   0.17045887919020208   0.25299833568389907   0.26524530532299945   0.13700938690197323   0.2718523081684915   0.38675974876899183   0.160389713713753   0.26086788834234115   0.6735764681619375   0.9189019833625843   0.3774269580722513   0.547222701963791   0.8545537250919473   0.6877260601676185   0.29072689717801514   0.6099100495020164   0.36843483206923866   0.21074576283830695   0.8320308078727779   0.5566129709438224   0.13402292179939068   0.6434379322467528   0.011694729906155166   0.9508038669108222   0.9635640426091886   0.3904395965628537   0.7464494245831557   0.8137944800088489   0.6917117344406971   0.0036798477938618877   0.5860597108694027   0.5529265916665078   0.018135266278759648   0.08477786443127755   0.20863275279715143   0.0057038897027167496
0.16358154118681242   0.39705180426365905   0.9179058556191363   0.3957938402007003   0.7951467091175738   0.18630604142535212   0.08587504774635829   0.8391808692568777   0.6611237873181831   0.5428681091785993   0.07418031784020312   0.8883770023460557   0.6975597447089945   0.1524285126157456   0.3277308932570474   0.0745825223372067   0.005848010268297324   0.14874866482188373   0.7416711823876447   0.5216559306706989   0.9877127439895377   0.0639708003906062   0.5330384295904933   0.5159520409679822   0.8241312028027252   0.6669189961269472   0.615132573971357   0.1201582007672819   0.028984493685151512   0.480612954701595   0.5292575262249987   0.2809773315104041   0.36786070636696844   0.9377448455229956   0.4550772083847956   0.39260032916434845   0.670300961657974   0.78531633290725   0.12734631512774816   0.31801780682714176   0.6644529513896766   0.6365676680853664   0.38567513274010345   0.7963618761564428   0.676740207400139   0.5725968676947601   0.8526367031496102   0.28040983518846063   0.8526090045974137   0.905677871567813   0.23750412917825317   0.16025163442117876   0.8236245109122622   0.425064916866218   0.7082466029532545   0.8792743029107747   0.45576380454529375   0.48732007134322236   0.2531693945684589   0.4866739737464262   0.7854628428873198   0.7020037384359723   0.12582307944071075   0.16865616691928442
0.12100989149764312   0.06543607035060597   0.7401479467006074   0.3722942907628416   0.4442696840975041   0.49283920265584585   0.8875112435509971   0.09188445557438092   0.5916606795000904   0.5871613310880328   0.6500071143727439   0.9316328211532021   0.7680361685878282   0.1620964142218148   0.9417605114194895   0.0523585182424275   0.31227236404253444   0.6747763428785924   0.6885911168510306   0.5656845444960014   0.5268095211552146   0.9727726044426201   0.5627680374103199   0.39702837757671694   0.40579962965757155   0.9073365340920142   0.8226200907097125   0.024734086813875344   0.9615299455600674   0.4144973314361684   0.9351088471587155   0.9328496312394944   0.369869266059977   0.8273360003481356   0.28510173278597145   0.0012168100862922754   0.6018330974721487   0.6652395861263207   0.343341221366482   0.9488582918438647   0.28956073342961436   0.9904632432477283   0.6547501045154513   0.38317374734786347   0.7627512122743997   0.017690638805108065   0.09198206710513154   0.9861453697711465   0.3569515826168282   0.11035410471309383   0.26936197639541903   0.9614112829572712   0.3954216370567608   0.6958567732769254   0.3342531292367036   0.028561651717776755   0.025552370996783806   0.8685207729287898   0.04915139645073216   0.027344841631484477   0.423719273524635   0.20328118680246912   0.7058101750842501   0.07848654978761971
0.13415854009502065   0.21281794355474085   0.05106007056879881   0.6953128024397562   0.3714073278206209   0.19512730474963277   0.9590780034636672   0.7091674326686097   0.014455745203792735   0.08477320003653896   0.6897160270682483   0.7477561497113385   0.619034108147032   0.3889164267596135   0.35546289783154467   0.7191944979935618   0.5934817371502481   0.5203956538308236   0.3063115013808125   0.6918496563620773   0.16976246362561312   0.31711446702835455   0.6005013262965623   0.6133631065744576   0.035603923530592475   0.10429652347361369   0.5494412557277635   0.9180503041347013   0.6641965957099716   0.9091692187239809   0.5903632522640962   0.2088828714660916   0.6497408505061788   0.824396018687442   0.900647225195848   0.46112672175475306   0.030706742359146874   0.4354795919278284   0.5451843273643033   0.7419322237611913   0.43722500520889873   0.9150839380970048   0.23887282598349083   0.05008256739911396   0.26746254158328564   0.5979694710686503   0.6383714996869285   0.43671946082465635   0.23185861805269314   0.49367294759503655   0.08893024395916507   0.5186691566899551   0.5676620223427216   0.5845037288710556   0.49856699169506885   0.30978628522386337   0.9179211718365428   0.7601077101836137   0.5979197664992209   0.8486595634691103   0.8872144294773959   0.32462811825578525   0.05273543913491759   0.10672733970791905
0.44998942426849714   0.40954418015878047   0.8138626131514267   0.05664477230880508   0.18252688268521153   0.8115747090901302   0.1754911134644982   0.6199253114841488   0.9506682646325184   0.31790176149509364   0.08656086950533314   0.10125615479419373   0.3830062422897968   0.733398032624038   0.5879938778102642   0.7914698695703304   0.46508507045325403   0.9732903224404243   0.9900741113110434   0.94281030610122   0.5778706409758582   0.6486622041846392   0.9373386721761258   0.8360829663933009   0.127881216707361   0.2391180240258587   0.12347605902469902   0.7794381940844959   0.9453543340221494   0.4275433149357285   0.9479849455602009   0.15951288260034718   0.994686069389631   0.10964155344063482   0.8614240760548677   0.05825672780615345   0.6116798270998343   0.3762435208165968   0.2734301982446034   0.2667868582358231   0.1465947566465802   0.40295319837617244   0.28335608693356007   0.3239765521346031   0.568724115670722   0.7542909941915333   0.3460174147574343   0.48789358574130215   0.44084289896336104   0.5151729701656746   0.22254135573273526   0.7084553916568063   0.49548856494121163   0.08762965522994619   0.27455641017253446   0.548942509056459   0.5008024955515806   0.9779881017893114   0.41313233411766676   0.4906857812503056   0.8891226684517464   0.6017445809727145   0.13970213587306338   0.2238989230144825
0.7425279118051662   0.19879138259654208   0.8563460489395033   0.8999223708798794   0.1738037961344441   0.4445003884050088   0.5103286341820691   0.41202878513857727   0.732960897171083   0.9293274182393341   0.28778727844933377   0.7035733934817711   0.23747233222987144   0.8416977630093879   0.013230868276799323   0.15463088442531198   0.7366698366782909   0.8637096612200765   0.6000985341591325   0.6639451031750063   0.8475471682265445   0.261965080247362   0.46039639828606915   0.4400461801605239   0.10501925642137834   0.06317369765081991   0.6040503493465659   0.5401238092806445   0.9312154602869342   0.6186733092458112   0.09372171516449682   0.12809502414206722   0.19825456311585118   0.689345891006477   0.8059344367151631   0.4245216306602962   0.9607822308859798   0.8476481279970891   0.7927035684383638   0.2698907462349842   0.2241123942076889   0.9839384667770126   0.19260503427923117   0.6059456430599778   0.3765652259811444   0.7219733865296506   0.732208635993162   0.16589946289945395   0.27154596955976606   0.6587996888788307   0.12815828664659612   0.6257756536188095   0.3403305092728318   0.04012637963301953   0.03443657148209931   0.49768062947674224   0.14207594615698063   0.3507804886265425   0.22850213476693626   0.0731589988164461   0.18129371527100088   0.5031323606294533   0.43579856632857256   0.803268252581462
0.957181321063312   0.5191938938524407   0.24319353204934138   0.1973226095214841   0.5806160950821676   0.7972205073227902   0.5109848960561794   0.03142314662203013   0.30907012552240154   0.13842081844395943   0.38282660940958324   0.40564749300322067   0.9687396162495697   0.09829443881093988   0.3483900379274839   0.9079668635264784   0.8266636700925891   0.7475139501843974   0.11988790316054766   0.8348078647100323   0.6453699548215882   0.2443815895549441   0.6840893368319751   0.03153961212857037   0.6881886337582762   0.7251876957025034   0.44089580478263374   0.8342170026070863   0.10757253867610861   0.9279671883797133   0.9299109087264543   0.8027938559850561   0.7985024131537071   0.7895463699357539   0.5470842993168711   0.39714636298183553   0.8297627969041373   0.691251931124814   0.1986942613893872   0.4891794994553571   0.00309912681154825   0.9437379809404166   0.07880635822883954   0.6543716347453249   0.35772917198996007   0.6993563913854725   0.39471702139686443   0.6228320226167545   0.6695405382316838   0.974168695682969   0.9538212166142307   0.7886150200096682   0.5619679995555753   0.046201507303255764   0.023910307887776306   0.9858211640246121   0.7634655864018682   0.2566551373675019   0.4768260085709052   0.5886748010427765   0.9337027894977309   0.5654032062426879   0.27813174718151795   0.09949530158741937
0.9306036626861827   0.6216652253022713   0.19932538895267843   0.44512366684209453   0.5728744906962225   0.9223088339167989   0.804608367555814   0.8222916442253401   0.9033339524645387   0.9481401382338298   0.8507871509415833   0.03367662421567188   0.34136595290896343   0.901938630930574   0.826876843053807   0.047855460191059865   0.5779003665070953   0.6452834935630721   0.35005083448290186   0.4591806591482834   0.6441975770093644   0.07988028732038427   0.07191908730138388   0.359685357560864   0.7135939143231818   0.4582150620181129   0.8725936983487055   0.9145616907187695   0.14071942362695924   0.535906228101314   0.06798533079289143   0.09227004649342939   0.23738547116242054   0.5877660898674842   0.2171981798513081   0.058593422277757504   0.896019518253457   0.6858274589369101   0.3903213367975011   0.01073796208669764   0.31811915174636185   0.040543965373837955   0.04027050231459923   0.5515573029384143   0.6739215747369974   0.9606636780534537   0.9683514150132153   0.1918719453775503   0.9603276604138157   0.5024486160353407   0.09575771666450991   0.27731025465878084   0.8196082367868565   0.9665423879340267   0.02777238587161847   0.18504020816535147   0.5822227656244359   0.37877629806654256   0.8105742060203104   0.12644678588759398   0.6862032473709788   0.6929488391296325   0.4202528692228093   0.11570882380089632
0.36808409562461697   0.6524048737557945   0.3799823669082101   0.564151520862482   0.6941625208876195   0.6917411957023407   0.4116309518949947   0.37227957548493174   0.7338348604738039   0.18929257966699997   0.31587323523048483   0.09496932082615088   0.9142266236869474   0.22275019173297325   0.2881008493588663   0.9099291126607995   0.33200385806251154   0.8439738936664307   0.477526643338556   0.7834823267732054   0.6458006106915327   0.15102505453679832   0.05727377411574668   0.6677735029723091   0.2777165150669158   0.49862018078100384   0.6772914072075367   0.10362198210982707   0.5835539941792963   0.8068789850786631   0.2656604553125419   0.7313424066248954   0.8497191337054925   0.6175864054116631   0.9497872200820571   0.6363730857987444   0.9354925100185449   0.3948362136786899   0.6616863707231908   0.7264439731379451   0.6034886519560334   0.5508623200122592   0.18415972738463482   0.9429616463647396   0.9576880412645007   0.39983726547546083   0.12688595326888813   0.2751881433924305   0.6799715261975848   0.9012170846944569   0.4495945460613515   0.17156616128260344   0.09641753201828858   0.09433809961579387   0.1839340907488096   0.44022375465770813   0.24669839831279616   0.4767516942041307   0.23414687066675247   0.8038506688589637   0.3112058882942512   0.08191548052544086   0.5724604999435617   0.07740669572101865
0.7077172363382178   0.5310531605131817   0.38830077255892687   0.13444504935627904   0.7500291950737171   0.13121589503772085   0.26141481929003874   0.8592569059638485   0.07005766887613224   0.22999881034326386   0.8118202732286872   0.6876907446812451   0.9736401368578437   0.13566071072747   0.6278861824798777   0.24746699002353703   0.7269417385450475   0.6589090165233392   0.3937393118131252   0.44361632116457334   0.4157358502507963   0.5769935359978984   0.8212788118695635   0.36620962544355473   0.7080186139125785   0.04594037548471668   0.4329780393106366   0.23176457608727566   0.9579894188388615   0.9147244804469958   0.17156322002059785   0.3725076701234271   0.8879317499627292   0.684725670103732   0.3597429467919106   0.684816925442182   0.9142916131048855   0.549064959376262   0.731856764312033   0.4373499354186449   0.187349874559838   0.8901559428529228   0.33811745249890773   0.9937336142540716   0.7716140243090417   0.3131624068550244   0.5168386406293443   0.6275239888105169   0.0635954103964632   0.2672220313703077   0.08386060131870762   0.3957594127232412   0.10560599155760178   0.35249755092331186   0.9122973812981098   0.02325174259981412   0.21767424159487261   0.6677718808195798   0.5525544345061992   0.33843481715763213   0.3033826284899871   0.11870692144331789   0.8206976701941663   0.9010848817389872
0.1160327539301491   0.22855097859039514   0.48258021769525855   0.9073512674849156   0.34441872962110737   0.9153885717353708   0.9657415770659143   0.2798272786743987   0.28082331922464415   0.648166540365063   0.8818809757472067   0.8840678659511575   0.1752173276670424   0.2956689894417512   0.9695835944490969   0.8608161233513434   0.9575430860721698   0.6278971086221713   0.41702915994289774   0.5223813061937113   0.6541604575821827   0.5091901871788534   0.5963314897487314   0.621296424454724   0.5381277036520336   0.2806392085884583   0.11375127205347292   0.7139451569698084   0.19370897403092618   0.36525063685308756   0.14800969498755862   0.4341178782954097   0.912885654806282   0.7170840964880245   0.266128719240352   0.5500500123442522   0.7376683271392396   0.42141510704627333   0.29654512479125505   0.6892338889929088   0.7801252410670698   0.793517998424102   0.8795159648483574   0.16685258279919754   0.12596478348488718   0.2843278112452486   0.28318447509962585   0.5455561583444735   0.5878370798328536   0.003688602656790265   0.16943320304615295   0.8316110013746651   0.3941281058019274   0.6384379658037027   0.02142350805859433   0.3974931230792554   0.4812424509956454   0.9213538693156782   0.7552947888182424   0.8474431107350032   0.7435741238564058   0.4999387622694049   0.45874966402698736   0.15820922174209445
0.9634488827893359   0.706420763845303   0.57923369917863   0.9913566389428969   0.8374840993044488   0.42209295260005436   0.29604922407900414   0.44580048059842337   0.24964701947159518   0.4184043499432641   0.12661602103285116   0.6141894792237582   0.8555189136696677   0.7799663841395613   0.10519251297425684   0.21669635614450286   0.3742764626740223   0.8586125148238831   0.34989772415601444   0.3692532454094996   0.6307023388176165   0.35867375255447825   0.8911480601290271   0.21104402366740518   0.6672534560282806   0.6522529887091754   0.3119143609503971   0.2196873847245083   0.8297693567238318   0.23016003610912097   0.015865136871392984   0.773886904126085   0.5801223372522366   0.8117556861658569   0.8892491158385418   0.15969742490232666   0.7246034235825689   0.03178930202629553   0.7840566028642849   0.9430010687578239   0.35032696090854654   0.17317678720241236   0.4341588787082705   0.5737478233483242   0.71962462209093   0.8145030346479342   0.5430108185792434   0.362703799680919   0.05237116606264941   0.1622500459387588   0.23109645762884629   0.14301641495641068   0.22260180933881762   0.9320900098296379   0.2152313207574533   0.36912951083032575   0.642479472086581   0.12033432366378093   0.3259822049189115   0.20943208592799908   0.9178760485040122   0.0885450216374854   0.5419256020546265   0.26643101717017525
0.5675490875954656   0.915368234435073   0.10776672334635601   0.6926831938218511   0.8479244655045356   0.1008651997871389   0.5647559047671126   0.32997939414093214   0.7955532994418862   0.9386151538483801   0.33365944713826634   0.18696297918452146   0.5729514901030686   0.006525144018742279   0.11842812638081306   0.8178334683541957   0.9304720180164876   0.8861908203549613   0.7924459214619016   0.6084013824261967   0.01259596951247547   0.797645798717476   0.25052031940727504   0.34197036525602137   0.44504688191700986   0.8822775642824029   0.14275359606091906   0.6492871714341703   0.5971224164124742   0.7814123644952641   0.5779976912938064   0.3193077772932381   0.8015691169705881   0.842797210646884   0.2443382441555401   0.1323447981087167   0.22861762686751944   0.8362720666281417   0.12591011777472705   0.314511329754521   0.2981456088510318   0.9500812462731804   0.3334641963128255   0.7061099473283243   0.28554963933855637   0.15243544755570435   0.08294387690555043   0.364139582072303   0.8405027574215465   0.2701578832733014   0.9401902808446314   0.7148524106381328   0.24338034100907224   0.48874551877803735   0.3621925895508249   0.39554463334489465   0.4418112240384842   0.6459483081311534   0.11785434539528482   0.26319983523617796   0.2131935971709648   0.8096762415030118   0.9919442276205578   0.948688505481657
0.915047988319933   0.8595949952298314   0.6584800313077322   0.2425785581533326   0.6294983489813766   0.7071595476741271   0.5755361544021819   0.8784389760810296   0.7889955915598301   0.4370016644008257   0.6353458735575505   0.16358656544289685   0.5456152505507579   0.9482561456227884   0.27315328400672556   0.7680419320980022   0.10380402651227365   0.3023078374916349   0.15529893861144076   0.5048420968618242   0.8906104293413089   0.49263159598862316   0.163354710990883   0.5561535913801673   0.9755624410213759   0.6330366007587916   0.5048746796831507   0.3135750332268347   0.34606409203999927   0.9258770530846646   0.9293385252809688   0.4351360571458051   0.5570685004801691   0.4888753886838389   0.2939926517234183   0.27154949170290826   0.011453249929411274   0.5406192430610506   0.02083936771669275   0.503507559604906   0.9076492234171376   0.23831140556941566   0.865540429105252   0.9986654627430818   0.017038794075828784   0.7456798095807925   0.702185718114369   0.4425118713629144   0.04147635305445291   0.11264320882200082   0.1973110384312183   0.1289368381360797   0.6954122610144536   0.18676615573733624   0.26797251315024945   0.6938007809902745   0.13834376053428452   0.6978907670534974   0.9739798614268311   0.4222512892873663   0.12689051060487322   0.1572715239924468   0.9531404937101384   0.9187437296824602
0.2192412871877356   0.9189601184230312   0.08760006460488638   0.9200782669393786   0.20220249311190683   0.1732803088422386   0.38541434649051737   0.4775663955764641   0.16072614005745392   0.0606371000202378   0.1881033080592991   0.3486295574403844   0.46531387904300026   0.8738709442829016   0.9201307949090496   0.6548287764501098   0.32697011850871577   0.1759801772294042   0.9461509334822186   0.23257748716274348   0.20007960790384252   0.018708653236957414   0.9930104397720801   0.31383375748028325   0.9808383207161069   0.09974853481392629   0.9054103751671938   0.3937554905409047   0.7786358276042001   0.9264682259716877   0.5199960286766764   0.9161890949644407   0.6179096875467462   0.8658311259514498   0.3318927206173773   0.5675595375240563   0.15259580850374596   0.9919601816685483   0.41176192570832765   0.9127307610739465   0.8256256899950302   0.8159800044391441   0.46561099222610913   0.680153273911203   0.6255460820911877   0.7972713512021867   0.472600552454029   0.36631951643091976   0.6447077613750807   0.6975228163882604   0.5671901772868352   0.972564025890015   0.8660719337708807   0.7710545904165728   0.04719414861015884   0.05637493092557438   0.2481622462241344   0.9052234644651229   0.7153014279927815   0.48881539340151814   0.09556643772038845   0.9132632827965745   0.3035395022844539   0.5760846323275717
0.26994074772535825   0.09728327835743047   0.8379285100583448   0.8959313584163687   0.6443946656341706   0.3000119271552438   0.36532795760431586   0.529611841985449   0.9996869042590899   0.6024891107669834   0.7981377803174806   0.557047816095434   0.13361497048820928   0.8314345203504107   0.7509436317073218   0.5006728851698595   0.8854527242640748   0.9262110558852877   0.03564220371454024   0.011857491768341449   0.7898862865436864   0.012947773088713182   0.7321027014300863   0.43577285944076977   0.5199455388183282   0.9156644947312828   0.8941741913717415   0.5398415010244011   0.8755508731841576   0.6156525675760389   0.5288462337674257   0.010229659038952144   0.8758639689250677   0.013163456809055552   0.7307084534499451   0.4531818429435182   0.7422489984368584   0.1817289364586449   0.9797648217426232   0.9525089577736586   0.8567962741727836   0.25551788057335717   0.944122618028083   0.9406514660053172   0.06690998762909711   0.242570107484644   0.21201991659799665   0.5048786065645474   0.546964448810769   0.3269056127533613   0.31784572522625515   0.9650371055401463   0.6714135756266114   0.7112530451773224   0.7889994914588295   0.9548074465011942   0.7955496067015437   0.6980895883682668   0.05829103800888452   0.5016256035576759   0.053300608264685266   0.5163606519096219   0.07852621626626131   0.5491166457840173
0.19650433409190174   0.2608427713362647   0.13440359823817835   0.6084651797787001   0.1295943464628046   0.018272663851620716   0.9223836816401817   0.10358657321415272   0.5826298976520357   0.6913670510982595   0.6045379564139265   0.13854946767400642   0.9112163220254242   0.9801140059209371   0.815538464955097   0.18374202117281227   0.11566671532388059   0.2820244175526703   0.7572474269462124   0.6821164176151363   0.062366107059195326   0.7656637656430484   0.6787212106799512   0.132999771831119   0.8658617729672936   0.5048209943067837   0.5443176124417728   0.5245345920524189   0.736267426504489   0.48654833045516305   0.6219339308015911   0.42094801883826616   0.15363752885245333   0.7951812793569035   0.017395974387664617   0.2823985511642597   0.24242120682702903   0.8150672734359665   0.20185750943256764   0.09865652999144746   0.12675449150314844   0.5330428558832961   0.4446100824863552   0.41654011237631117   0.06438838444395312   0.7673790902402478   0.7658888718064041   0.2835403405451921   0.1985266114766595   0.262558095933464   0.2215712593646313   0.7590057484927732   0.4622591849721705   0.7760097654783009   0.5996373285630402   0.3380577296545071   0.3086216561197172   0.9808284861213974   0.5822413541753756   0.05565917849024738   0.06620044929268815   0.1657612126854309   0.3803838447428079   0.9570026484987999
0.9394459577895397   0.6327183568021347   0.9357737622564527   0.5404625361224887   0.8750575733455866   0.865339266561887   0.16988489045004862   0.2569221955772966   0.676530961868927   0.602781170628423   0.9483136310854173   0.4979164470845234   0.21427177689675656   0.826771405150122   0.34867630252237714   0.15985871743001626   0.9056501207770393   0.8459429190287246   0.7664349483470015   0.10419953893976888   0.8394496714843512   0.6801817063432938   0.3860511036041937   0.14719689044096895   0.9000037136948115   0.047463349541159   0.450277341347741   0.6067343543184802   0.02494614034922493   0.182124082979272   0.2803924508976923   0.34981215874118354   0.34841517848029785   0.579342912350849   0.332078819812275   0.8518957116566602   0.13414340158354127   0.752571507200727   0.9834025172898979   0.6920369942266439   0.2284932808065019   0.9066285881720023   0.21696756894289626   0.587837455286875   0.38904360932215065   0.22644688182870856   0.8309164653387026   0.4406405648459061   0.4890398956273392   0.17898353228754954   0.3806391239909616   0.8339062105274259   0.46409375527811425   0.9968594493082775   0.10024667309326926   0.4840940517862423   0.11567857679781639   0.4175165369574286   0.7681678532809942   0.6321983401295822   0.9815351752142751   0.6649450297567017   0.7847653359910964   0.9401613459029382
0.7530418944077732   0.7583164415846994   0.5677977670482002   0.3523238906160632   0.36399828508562254   0.5318695597559908   0.7368813017094975   0.9116833257701571   0.8749583894582834   0.3528860274684413   0.35624217771853595   0.07777711524273119   0.41086463418016916   0.3560265781601637   0.25599550462526666   0.5936830634564888   0.29518605738235276   0.9385100412027351   0.4878276513442724   0.9614847233269067   0.3136508821680776   0.27356501144603346   0.703062315353176   0.021323377423968472   0.5606089877603044   0.5152485698613342   0.1352645483049759   0.6689994868079053   0.19661070267468192   0.9833790101053433   0.39838324659547836   0.7573161610377482   0.32165231321639853   0.630492982636902   0.04214106887694242   0.679539045795017   0.9107876790362294   0.27446640447673837   0.7861455642516758   0.08585598233852815   0.6156016216538767   0.33595636327400324   0.2983179129074034   0.12437125901162145   0.30195073948579904   0.06239135182796976   0.5952555975542274   0.10304788158765298   0.7413417517254945   0.5471427819666357   0.4599910492492515   0.43404839477974766   0.5447310490508126   0.5637637718612923   0.06160780265377315   0.6767322337419995   0.2230787358344141   0.9332707892243903   0.01946673377683073   0.9971931879469825   0.3122910567981847   0.6588043847476519   0.23332116952515497   0.9113372056084543
0.696689435144308   0.3228480214736487   0.9350032566177516   0.7869659465968329   0.394738695658509   0.26045666964567893   0.3397476590635242   0.68391806500918   0.6533969439330144   0.7133138876790432   0.8797566098142727   0.24986967022943224   0.10866589488220178   0.14955011581775096   0.8181488071604995   0.5731374364874328   0.8855871590477877   0.21627932659336066   0.7986820733836688   0.5759442485404502   0.573296102249603   0.5574749418457088   0.5653609038585139   0.6646070429319959   0.876606667105295   0.23462692037206   0.6303576472407623   0.8776410963351631   0.481867971446786   0.9741702507263811   0.2906099881772381   0.19372303132598312   0.8284710275137716   0.2608563630473378   0.4108533783629653   0.9438533610965509   0.7198051326315698   0.11130624722958682   0.5927045712024658   0.3707159246091181   0.8342179735837821   0.8950269206362261   0.7940224978187969   0.7947716760686678   0.2609218713341791   0.3375519787905174   0.228661593960283   0.13016463313667193   0.3843152042288841   0.1029250584184574   0.5983039467195207   0.2525235368015089   0.902447232782098   0.1287548076920763   0.3076939585422826   0.05880050547552578   0.07397620526832652   0.8678984446447385   0.8968405801793172   0.11494714437897491   0.35417107263675673   0.7565921974151517   0.30413600897685156   0.7442312197698567
0.5199530990529746   0.8615652767789256   0.5101135111580546   0.9494595437011889   0.25903122771879555   0.5240132979884081   0.28145191719777163   0.819294910564517   0.8747160234899115   0.42108823956995073   0.6831479704782509   0.566771373763008   0.9722687907078135   0.2923334318778744   0.37545401193596833   0.5079708682874823   0.8982925854394869   0.4244349872331359   0.47861343175665105   0.39302372390850737   0.5441215128027301   0.6678427898179842   0.17447742277979952   0.6487925041386506   0.024168413749755514   0.8062775130390586   0.6643639116217449   0.6993329604374617   0.7651371860309599   0.28226421505065047   0.3829119944239732   0.8800380498729448   0.8904211625410484   0.8611759754806997   0.6997640239457222   0.3132666761099367   0.9181523718332351   0.5688425436028253   0.32431001200975396   0.8052958078224544   0.01985978639374814   0.1444075563696894   0.8456965802531029   0.412272083913947   0.475738273591018   0.47656476655170527   0.6712191574733033   0.7634795797752963   0.45156985984126247   0.6702872535126466   0.006855245851558443   0.06414661933783469   0.6864326738103025   0.3880230384619962   0.6239432514275852   0.18410856946488996   0.7960115112692541   0.5268470629812965   0.9241792274818629   0.8708418933549533   0.877859139436019   0.9580045193784712   0.599869215472109   0.0655460855324989
0.8579993530422709   0.8135969630087818   0.7541726352190061   0.6532740016185519   0.3822610794512529   0.3370321964570765   0.0829534777457028   0.8897944218432555   0.9306912196099905   0.6667449429444299   0.07609823189414436   0.8256478025054208   0.24425854579968795   0.27872190448243367   0.45215498046655916   0.6415392330405308   0.44824703453043385   0.7518748415011371   0.5279757529846962   0.7706973396855775   0.5703878950944149   0.793870322122666   0.9281065375125872   0.7051512541530787   0.712388542052144   0.9802733591138842   0.1739339022935811   0.05187725253452678   0.33012746260089104   0.6432411626568076   0.09098042454787829   0.1620828306912713   0.3994362429909006   0.9764962197123779   0.014882192653733941   0.3364350281858505   0.15517769719121266   0.6977743152299442   0.5627272121871748   0.6948957951453197   0.7069306626607788   0.945899473728807   0.03475145920247857   0.9241984554597421   0.13654276756636394   0.152029151606141   0.10664492168989134   0.21904720130666347   0.42415422551422   0.17175579249225678   0.9327110193963103   0.1671699487721367   0.09402676291332894   0.5285146298354491   0.8417305948484319   0.005087118080865388   0.6945905199224284   0.5520184101230713   0.826848402194698   0.6686520898950149   0.5394128227312157   0.8542440948931271   0.2641211900075232   0.9737562947496952
0.832482160070437   0.9083446211643201   0.22936973080504466   0.049557839289953054   0.695939392504073   0.7563154695581791   0.12272480911515331   0.8305106379832896   0.271785166989853   0.5845596770659223   0.19001378971884306   0.6633406892111529   0.17775840407652407   0.05604504723047319   0.3482831948704111   0.6582535711302875   0.48316788415409573   0.5040266371074019   0.5214347926757131   0.9896014812352726   0.94375506142288   0.6497825422142748   0.25731360266818987   0.01584518648557744   0.1112729013524431   0.7414379210499548   0.027943871863145203   0.9662873471956244   0.4153335088483701   0.9851224514917757   0.9052190627479919   0.1357767092123348   0.14354834185851711   0.40056277442585336   0.7152052730291488   0.4724360200011819   0.9657899377819931   0.34451772719538015   0.36692207815873773   0.8141824488708944   0.48262205362789734   0.8404910900879783   0.8454872854830247   0.8245809676356218   0.5388669922050173   0.19070854787370342   0.5881736828148348   0.8087357811500444   0.4275940908525742   0.4492706268237487   0.5602298109516896   0.8424484339544199   0.01226058200420409   0.464148175331973   0.6550107482036978   0.7066717247420852   0.8687122401456869   0.06358540090611965   0.9398054751745488   0.23423570474090324   0.902922302363694   0.7190676737107394   0.5728833970158111   0.4200532558700088
0.4203002487357966   0.8785765836227613   0.7273961115327865   0.595472288234387   0.8814332565307793   0.6878680357490579   0.13922242871795168   0.7867365070843426   0.4538391656782051   0.23859740892530917   0.5789926177662621   0.9442880731299227   0.441578583674001   0.7744492335933362   0.9239818695625643   0.2376163483878375   0.572866343528314   0.7108638326872165   0.9841763943880155   0.0033806436469342683   0.66994404116462   0.991796158976477   0.41129299737220437   0.5833273877769255   0.24964379242882348   0.11321957535371577   0.6838968858394179   0.9878550995425385   0.3682105358980442   0.42535153960465794   0.5446744571214662   0.20111859245819583   0.9143713702198392   0.18675413067934876   0.9656818393552041   0.25683051932827317   0.4727927865458382   0.41230489708601264   0.0416999697926398   0.019214170940435656   0.8999264430175241   0.7014410643987962   0.057523575404624286   0.01583352729350139   0.22998240185290406   0.7096449054223191   0.6462305780324199   0.4325061395165759   0.9803386094240806   0.5964253300686033   0.962333692193002   0.4446510399740375   0.6121280735260364   0.1710737904639454   0.41765923507153574   0.24353244751584163   0.6977567033061972   0.9843196597845967   0.45197739571633155   0.9867019281875685   0.22496391676035907   0.572014762698584   0.41027742592369176   0.9674877572471329
0.3250374737428349   0.8705736982997879   0.3527538505190675   0.9516542299536315   0.09505507188993084   0.16092879287746875   0.7065232724866476   0.5191480904370555   0.11471646246585027   0.5645034628088654   0.7441895802936456   0.07449705046301805   0.502588388939814   0.39342967234492005   0.32653034522210983   0.8309646029471764   0.8048316856336167   0.40911001256032337   0.8745529495057782   0.8442626747596079   0.5798677688732576   0.8370952498617393   0.4642755235820865   0.8767749175124752   0.2548302951304227   0.9665215515619515   0.11152167306301901   0.9251206875588437   0.1597752232404919   0.8055927586844828   0.40499840057637143   0.4059725971217882   0.04505876077464162   0.2410892958756173   0.6608088202827258   0.3314755466587701   0.5424703718348277   0.8476596235306973   0.334278475060616   0.5005109437115938   0.737638686201211   0.4385496109703739   0.4597255255548377   0.6562482689519857   0.15777091732795337   0.6014543611086345   0.9954500019727512   0.7794733514395107   0.9029406221975307   0.634932809546683   0.8839283289097322   0.854352663880667   0.7431653989570387   0.8293400508622003   0.4789299283333608   0.4483800667588788   0.6981066381823972   0.588250754986583   0.818121108050635   0.11690452010010871   0.1556362663475694   0.7405911314558856   0.483842632990019   0.616393576388515
0.4179975801463584   0.30204152048551175   0.024117107435181317   0.9601453074365293   0.26022666281840506   0.7005871593768772   0.028667105462430127   0.18067195599701852   0.3572860406208744   0.06565434983019422   0.14473877655269793   0.3263192921163515   0.6141206416638356   0.23631429896799394   0.6658088482193372   0.8779392253574727   0.9160140034814385   0.648063543981411   0.8476877401687022   0.7610347052573639   0.7603777371338691   0.9074724125255254   0.3638451071786832   0.14464112886884897   0.3423801569875107   0.6054308920400135   0.3397279997435019   0.18449582143231977   0.08215349416910564   0.9048437326631363   0.31106089428107175   0.0038238654353012404   0.7248674535482312   0.8391893828329421   0.16632211772837383   0.6775045733189498   0.11074681188439559   0.6028750838649481   0.5005132695090366   0.799565347961477   0.19473280840295706   0.9548115398835372   0.6528255293403344   0.038530642704113056   0.43435507126908796   0.047339127358011865   0.28898042216165126   0.893889513835264   0.0919749142815773   0.4419082353179983   0.9492524224181493   0.7093936924029443   0.009821420112471661   0.5370645026548619   0.6381915281370776   0.705569826967643   0.28495396656424044   0.6978751198219199   0.4718694104087038   0.02806525364869335   0.17420715467984485   0.09500003595697168   0.9713561408996672   0.22849990568721631
0.9794743462768878   0.1401884960734345   0.31853061155933265   0.18996926298310327   0.5451192750077998   0.09284936871542263   0.029550189397681413   0.2960797491478392   0.4531443607262225   0.6509411333974243   0.08029776697953206   0.5866860567448949   0.4433229406137508   0.11387663074256235   0.4421062388424545   0.8811162297772518   0.15836897404951042   0.4160015109206425   0.9702368284337507   0.8530509761285585   0.9841618193696656   0.3210014749636708   0.9988806875340835   0.6245510704413422   0.004687473092777795   0.18081297889023634   0.680350075974751   0.4345818074582389   0.459568198084978   0.0879636101748137   0.6507998865770696   0.1385020583103997   0.006423837358755473   0.43702247677738937   0.5705021195975375   0.5518160015655048   0.5631008967450046   0.32314584603482704   0.128395880755083   0.670699771788253   0.4047319226954942   0.9071443351141846   0.1581590523213323   0.8176487956596945   0.4205701033258286   0.5861428601505138   0.15927836478724872   0.19309772521835236   0.41588263023305083   0.40532988126027736   0.47892828881249777   0.7585159177601135   0.9563144321480729   0.31736627108546367   0.8281284022354283   0.6200138594497138   0.9498905947893174   0.8803437943080743   0.2576262826378908   0.06819785788420901   0.38678969804431274   0.5571979482732472   0.1292304018828078   0.39749808609595605
0.9820577753488186   0.6500536131590627   0.9710713495614756   0.5798492904362615   0.5614876720229899   0.06391075300854902   0.8117929847742268   0.38675156521790915   0.1456050417899391   0.6585808717482716   0.332864695961729   0.6282356474577957   0.18929060964186625   0.341214600662808   0.5047362937263008   0.008221788008081833   0.2394000148525489   0.4608708063547337   0.24711001108840996   0.9400239301238729   0.8526103168082362   0.9036728580814865   0.11787960920560214   0.5425258440279168   0.8705525414594176   0.2536192449224237   0.14680825964412664   0.9626765535916553   0.3090648694364277   0.1897084919138747   0.33501527486989985   0.5759249883737462   0.16345982764648856   0.5311276201656031   0.0021505789081708287   0.9476893409159505   0.9741692180046223   0.18991301950279507   0.4974142851818701   0.9394675529078687   0.7347692031520734   0.7290422131480614   0.2503042740934601   0.9994436227839958   0.8821588863438373   0.8253693550665749   0.13242466488785798   0.45691777875607903   0.011606344884419677   0.5717501101441512   0.9856164052437313   0.49424122516442376   0.7025414754479921   0.3820416182302765   0.6506011303738315   0.9183162367906776   0.5390816478015035   0.8509139980646734   0.6484505514656607   0.9706268958747272   0.5649124297968812   0.6610009785618783   0.15103626628379058   0.031159342966858496
0.8301432266448077   0.931958765413817   0.9007319921903305   0.031715720182862665   0.9479843403009705   0.10658941034724208   0.7683073273024725   0.5747979414267836   0.9363779954165508   0.5348393002030909   0.7826909220587411   0.08055671626235986   0.23383651996855875   0.1527976819728144   0.13208979168490967   0.16224047947168221   0.6947548721670553   0.30188368390814097   0.48363924021924903   0.19161358359695507   0.12984244237017417   0.6408827053462626   0.3326029739354584   0.16045424063009656   0.29969921572536645   0.7089239399324456   0.43187098174512795   0.1287385204472339   0.351714875424396   0.6023345295852035   0.6635636544426555   0.5539405790204502   0.41533688000784524   0.06749522938211264   0.8808727323839143   0.4733838627580904   0.18150036003928652   0.9146975474092982   0.7487829406990046   0.3111433832864082   0.4867454878722312   0.6128138635011573   0.26514370047975566   0.11952979968945315   0.35690304550205704   0.9719311581548946   0.9325407265442972   0.9590755590593566   0.05720382977669054   0.26300721822244905   0.5006697447991693   0.8303370386121227   0.7054889543522945   0.6606726886372455   0.8371060903565137   0.2763964595916724   0.2901520743444493   0.5931774592551329   0.9562333579725995   0.803012596833582   0.10865171430516275   0.6784799118458347   0.2074504172735948   0.4918692135471738
0.6219062264329316   0.06566604834467737   0.9423067167938391   0.3723394138577206   0.26500318093087455   0.09373489018978272   0.009765990249541964   0.413263854798364   0.207799351154184   0.8307276719673337   0.5090962454503727   0.5829268161862413   0.5023103968018895   0.17005498333008814   0.671990155093859   0.3065303565945689   0.21215832245744023   0.5768775240749553   0.7157567971212595   0.5035177597609869   0.10350660815227747   0.8983976122291206   0.5083063798476647   0.011648546213813178   0.4816003817193459   0.8327315638844432   0.5659996630538254   0.6393091323560925   0.21659720078847136   0.7389966736946606   0.5562336728042835   0.22604527755772857   0.008797849634287347   0.9082690017273268   0.0471374273539108   0.6431184613714872   0.5064874528323978   0.7382140183972388   0.37514727226005185   0.3365881047769183   0.2943291303749576   0.16133649432228345   0.6593904751387923   0.8330703450159314   0.19082252222268017   0.2629388820931628   0.15108409529112773   0.8214217988021182   0.7092221405033343   0.43020731820871955   0.5850844322373022   0.18211266644602564   0.49262493971486293   0.691210644514059   0.02885075943301876   0.9560673888882971   0.48382709008057556   0.7829416427867322   0.9817133320791079   0.3129489275168098   0.9773396372481777   0.0447276243894934   0.6065660598190561   0.9763608227398914
0.6830105068732201   0.8833911300672099   0.9471755846802637   0.14329047772396009   0.4921879846505399   0.6204522479740472   0.796091489389136   0.3218686789218419   0.7829658441472056   0.19024492976532761   0.21100705715183368   0.13975601247581623   0.29034090443234273   0.49903428525126864   0.18215629771881492   0.18368862358751917   0.8065138143517672   0.7160926424645365   0.20044296563970695   0.8707396960707093   0.8291741771035894   0.6713650180750431   0.5938769058206509   0.8943788733308179   0.14616367023036936   0.7879738880078331   0.6467013211403871   0.7510883956068578   0.6539756855798294   0.16752164003378597   0.8506098317512512   0.42921971668501585   0.8710098414326238   0.9772767102684583   0.6396027745994175   0.28946370420919965   0.5806689370002811   0.4782424250171897   0.4574464768806026   0.10577508062168048   0.7741551226485139   0.7621497825526532   0.25700351124089565   0.23503538455097114   0.9449809455449245   0.09078476447761015   0.6631266054202448   0.3406565112201533   0.7988172753145552   0.30281087646977706   0.016425284279857618   0.5895681156132956   0.14484158973472572   0.13528923643599106   0.1658154525286064   0.16034839892827968   0.2738317483021019   0.15801252616753272   0.5262126779291889   0.87088469471908   0.6931628113018208   0.679770101150343   0.06876620104858627   0.7651096140973995
0.9190076886533067   0.9176203185976898   0.8117626898076906   0.5300742295464285   0.9740267431083822   0.8268355541200796   0.14863608438744585   0.18941771832627513   0.17520946779382698   0.5240246776503026   0.13221080010758823   0.5998496027129796   0.030367878059101287   0.3887354412143115   0.9663953475789818   0.4395012037846999   0.7565361297569995   0.23072291504677878   0.4401826696497929   0.5686165090656199   0.0633733184551787   0.5509528138964358   0.37141646860120664   0.8035068949682204   0.14436562980187195   0.633332495298746   0.5596537787935161   0.2734326654217919   0.1703388866934898   0.8064969411786664   0.41101769440607017   0.0840149470955168   0.9951294188996628   0.28247226352836385   0.27880689429848193   0.4841653443825372   0.9647615408405615   0.8937368223140524   0.3124115467195001   0.04466414059783731   0.20822541108356207   0.6630139072672736   0.8722288770697072   0.47604763153221746   0.14485209262838336   0.11206109337083782   0.5008124084685005   0.6725407365639972   0.0004864628265114064   0.4787285980720918   0.9411586296749845   0.3991080711422052   0.8301475761330216   0.6722316568934253   0.5301409352689144   0.31509312404668843   0.8350181572333588   0.3897593933650615   0.2513340409704324   0.8309277796641512   0.8702566163927973   0.4960225710510091   0.9389224942509322   0.7862636390663139
0.6620312053092352   0.8330086637837355   0.06669361718122507   0.31021600753409645   0.5171791126808519   0.7209475704128977   0.5658812087127245   0.6376752709700994   0.5166926498543405   0.2422189723408059   0.6247225790377401   0.23856719982789412   0.6865450737213189   0.5699873154473806   0.09458164376882572   0.9234740757812057   0.85152691648796   0.18022792208231905   0.8432476027983933   0.09254629611705449   0.9812703000951627   0.68420535103131   0.9043251085474611   0.3062826570507406   0.31923909478592744   0.8511966872475745   0.837631491366236   0.9960666495166441   0.8020599821050756   0.13024911683467671   0.2717502826535115   0.35839137854654485   0.2853673322507351   0.8880301444938709   0.6470277036157714   0.11982417871865071   0.5988222585294163   0.3180428290464903   0.5524460598469457   0.196350102937445   0.7472953420414562   0.13781490696417126   0.7091984570485523   0.10380380682039053   0.7660250419462935   0.45360955593286134   0.8048733485010913   0.7975211497696499   0.44678594716036607   0.6024128686852869   0.9672418571348553   0.8014545002530058   0.6447259650552906   0.4721637518506102   0.6954915744813438   0.44306312170646095   0.35935863280455543   0.5841336073567394   0.048463870865572384   0.3232389429878102   0.7605363742751392   0.2660907783102491   0.4960178110186267   0.1268888400503652
0.013241032233682965   0.12827587134607782   0.7868193539700743   0.023085033229974662   0.24721599028738944   0.6746663154132165   0.981946005468983   0.22556388346032474   0.8004300431270234   0.07225344672792959   0.014704148334127719   0.424109383207319   0.15570407807173284   0.6000896948773194   0.3192125738527839   0.981046261500858   0.7963454452671774   0.015956087520580038   0.27074870298721154   0.6578073185130479   0.03580907099203825   0.749865309210331   0.7747308919685848   0.5309184784626826   0.022568038758355283   0.6215894378642531   0.9879115379985105   0.507833445232708   0.7753520484709658   0.9469231224510366   0.005965532529527544   0.2822695617723832   0.9749220053439425   0.874669675723107   0.9912613841953998   0.8581601785650642   0.8192179272722097   0.27457998084578766   0.6720488103426159   0.8771139170642062   0.022872482005032193   0.25862389332520763   0.4013001073554044   0.2193065985511584   0.987063411012994   0.5087585841148766   0.6265692153868195   0.6883881200884757   0.9644953722546387   0.8871691462506235   0.638657677388309   0.18055467485576776   0.18914332378367282   0.9402460237995869   0.6326921448587814   0.8982851130833845   0.21422131843973036   0.06557634807647979   0.6414307606633817   0.04012493451832028   0.3950033911675207   0.7909963672306921   0.9693819503207657   0.16301101745411406
0.37213090916248853   0.5323724739054845   0.5680818429653613   0.9437044189029556   0.3850674981494946   0.023613889790607825   0.9415126275785417   0.2553162988144799   0.42057212589485593   0.13644474353998431   0.30285495019023273   0.07476162395871216   0.2314288021111831   0.19619871974039746   0.6701628053314512   0.17647651087532762   0.017207483671452747   0.13062237166391766   0.028732044668069626   0.13635157635700734   0.622204092503932   0.33962600443322555   0.05935009434730391   0.9733405589028933   0.2500731833414435   0.8072535305277411   0.4912682513819426   0.02963613999993761   0.8650056851919489   0.7836396407371332   0.5497556238034008   0.7743198411854577   0.444433559297093   0.647194897197149   0.2469006736131681   0.6995582172267455   0.2130047571859099   0.45099617745675147   0.5767378682817168   0.5230817063514179   0.19579727351445714   0.3203738057928338   0.5480058236136471   0.38673012999441053   0.5735931810105251   0.9807478013596083   0.48865572926634326   0.41338957109151725   0.3235199976690816   0.1734942708318672   0.9973874778844007   0.3837534310915796   0.4585143124771327   0.3898546300947339   0.44763185408099987   0.609433589906122   0.014080753180039741   0.742659732897585   0.20073118046783178   0.9098753726793765   0.8010759959941298   0.29166355544083356   0.623993312186115   0.38679366632795853
0.6052787224796727   0.9712897496479997   0.07598748857246777   0.00006353633354803478   0.03168554146914759   0.9905419482883915   0.5873317593061245   0.5866739652420309   0.7081655438000659   0.8170476774565243   0.5899442814217238   0.2029205341504512   0.24965123132293324   0.42719304736179037   0.1423124273407239   0.5934869442443292   0.2355704781428935   0.6845333144642054   0.9415812468728921   0.6836115715649528   0.4344944821487636   0.3928697590233718   0.31758793468677715   0.29681790523699425   0.8292157596690909   0.42158000937537204   0.2416004461143094   0.29675436890344625   0.7975302181999433   0.43103806108698056   0.654268686808185   0.7100804036614154   0.08936467439987737   0.6139903836304562   0.06432440538646113   0.5071598695109643   0.8397134430769442   0.18679733626866588   0.9220119780457372   0.913672925266635   0.6041429649340506   0.5022640218044605   0.9804307311728451   0.23006135370168215   0.16964848278528702   0.1093942627810887   0.6628427964860679   0.9332434484646879   0.3404327231161961   0.6878142534057167   0.4212423503717585   0.6364890795612417   0.5429025049162527   0.25677619231873605   0.7669736635635735   0.9264086758998262   0.45353783051637536   0.6427858086882798   0.7026492581771124   0.419248806388862   0.6138243874394312   0.45598847241961393   0.7806372801313752   0.5055758811222271
0.00968142250538057   0.9537244506151534   0.8002065489585302   0.2755145274205449   0.8400329397200935   0.8443301878340648   0.13736375247246224   0.34227107895585696   0.4996002166038975   0.1565159344283481   0.7161214021007037   0.7057819993946153   0.9566977116876447   0.899739742109612   0.9491477385371301   0.779373323494789   0.5031598811712693   0.2569539334213322   0.24649848036001767   0.360124517105927   0.8893354937318382   0.8009654610017183   0.4658612002286424   0.8545486359837   0.8796540712264576   0.8472410103865649   0.6656546512701123   0.5790341085631551   0.03962113150636401   0.0029108225525001073   0.52829089879765   0.23676302960729811   0.5400209149024665   0.846394888124152   0.8121694966969463   0.5309810302126828   0.5833232032148218   0.94665514601454   0.8630217581598162   0.7516077067178938   0.08016332204355245   0.6897012125932078   0.6165232777997985   0.39148318961196676   0.19082782831171433   0.8887357515914895   0.15066207757115607   0.5369345536282668   0.31117375708525674   0.04149474120492468   0.4850074263010438   0.9579004450651116   0.27155262557889276   0.038583918652424574   0.9567165275033938   0.7211374154578135   0.7315317106764262   0.19218903052827255   0.14454703080644746   0.19015638524513073   0.1482085074616044   0.24553388451373256   0.28152527264663124   0.43854867852723695
0.06804518541805195   0.5558326719205248   0.6650019948468328   0.04706548891527021   0.8772173571063376   0.6670969203290352   0.5143399172756767   0.5101309352870035   0.5660436000210809   0.6256021791241106   0.029332490974632898   0.5522304902218917   0.29449097444218814   0.587018260471686   0.07261596347123914   0.8310930747640782   0.5629592637657619   0.39482922994341346   0.9280689326647917   0.6409366895189474   0.41475075630415753   0.1492953454296809   0.6465436600181604   0.20238801099171055   0.34670557088610554   0.593462673509156   0.9815416651713277   0.15532252207644034   0.46948821377976796   0.9263657531801208   0.467201747895651   0.6451915867894369   0.9034446137586871   0.30076357405601023   0.4378692569210181   0.09296109656754513   0.6089536393164989   0.7137453135843242   0.3652532934497789   0.2618680218034669   0.04599437555073705   0.31891608364091073   0.43718436078498724   0.6209313322845194   0.6312436192465796   0.16962073821122986   0.7906407007668268   0.41854332129280886   0.28453804836047397   0.5761580647020738   0.8090990355954991   0.26322079921636854   0.815049834580706   0.6497923115219529   0.3418972876998482   0.6180292124269317   0.911605220822019   0.3490287374659427   0.9040280307788301   0.5250681158593865   0.30265158150552   0.6352834238816185   0.5387747373290511   0.2632000940559196
0.256657205954783   0.3163673402407078   0.10159037654406393   0.6422687617714001   0.6254135867082035   0.1467466020294779   0.31094967577723714   0.22372544047859133   0.34087553834772943   0.5705885373274041   0.501850640181738   0.9605046412622228   0.5258257037670234   0.9207962258054512   0.1599533524818898   0.3424754288352912   0.6142204829450044   0.5717674883395084   0.2559253217030597   0.8174073129759047   0.3115689014394844   0.9364840644578899   0.7171505843740086   0.5542072189199851   0.05491169548470144   0.6201167242171821   0.6155602078299446   0.9119384571485849   0.429498108776498   0.47337012218770425   0.3046105320527075   0.6882130166699936   0.0886225704287686   0.9027815848603001   0.8027598918709695   0.7277083754077708   0.5627968666617452   0.981985359054849   0.6428065393890797   0.38523294657247964   0.9485763837167408   0.41021787071534055   0.38688121768601996   0.5678256335965749   0.6370074822772565   0.4737338062574506   0.6697306333120114   0.013618414676589821   0.5820957867925549   0.8536170820402684   0.05417042548206682   0.10167995752800489   0.15259767801605695   0.3802469598525642   0.7495598934293594   0.4134669408580113   0.06397510758728833   0.47746537499226405   0.9468000015583898   0.6857585654502405   0.5011782409255431   0.49548001593741503   0.3039934621693101   0.30052561887776086
0.5526018572088023   0.0852621452220745   0.9171122444832901   0.732699985281186   0.9155943749315459   0.6115283389646239   0.2473816111712787   0.7190815706045961   0.3334985881389909   0.7579112569243555   0.1932111856892119   0.6174016130765912   0.180900910122934   0.3776642970717912   0.44365129225985256   0.20393467221857992   0.11692580253564566   0.9001989220795272   0.4968512907014627   0.5181761067683395   0.6157475616101026   0.40471890614211214   0.19285782853215264   0.21765048789057861   0.06314570440130025   0.31945676092003766   0.2757455840488625   0.4849505026093927   0.14755132946975436   0.7079284219554138   0.028363972877583805   0.7658689320047967   0.8140527413307634   0.9500171650310584   0.8351527871883719   0.14846731892820542   0.6331518312078295   0.5723528679592671   0.3915014949285194   0.9445326467096256   0.5162260286721837   0.6721539458797399   0.8946502042270567   0.4263565399412861   0.9004784670620812   0.2674350397376278   0.701792375694904   0.20870605205070744   0.8373327626607809   0.9479782788175901   0.4260467916460415   0.7237555494413147   0.6897814331910266   0.2400498568621763   0.3976828187684577   0.9578866174365182   0.8757286918602631   0.29003269183111796   0.5625300315800857   0.8094192985083127   0.24257686065243378   0.7176798238718508   0.1710285366515664   0.8648866517986872
0.72635083198025   0.04552587799211092   0.27637833242450977   0.43853011185740115   0.8258723649181688   0.7780908382544831   0.5745859567296058   0.2298240598066937   0.9885396022573879   0.8301125594368931   0.14853916508356424   0.5060685103653789   0.29875816906636127   0.5900627025747167   0.7508563463151066   0.5481818929288608   0.42302947720609807   0.3000300107435988   0.1883263147350208   0.7387625944205481   0.1804526165536643   0.582350186871748   0.017297778083454403   0.8738759426218609   0.45410178457341427   0.5368243088796371   0.7409194456589446   0.43534583076445976   0.6282294196552455   0.7587334706251538   0.16633348892933889   0.20552177095776605   0.6396898173978576   0.9286209111882608   0.01779432384577464   0.6994532605923871   0.34093164833149636   0.3385582086135441   0.26693797753066806   0.15127136766352625   0.9179021711253983   0.03852819786994526   0.07861166279564728   0.41250877324297813   0.737449554571734   0.4561780109981973   0.06131388471219288   0.5386328306211172   0.28334776999831973   0.9193537021185603   0.3203944390532482   0.10328699985665751   0.6551183503430742   0.1606202314934064   0.15406095012390936   0.8977652288988914   0.015428532945216612   0.2319993203051456   0.1362666262781347   0.19831196830650438   0.6744968846137203   0.8934411116916016   0.8693286487474666   0.047040600642978124
0.756594713488322   0.8549129138216562   0.7907169859518194   0.6345318273999999   0.019145158916587916   0.39873490282345897   0.7294031012396265   0.09589899677888271   0.7357973889182682   0.4793812007048987   0.4090086621863782   0.9926119969222252   0.08067903857519396   0.3187609692114923   0.25494771206246886   0.09484676802333371   0.06525050562997735   0.08676164890634669   0.11868108578433417   0.8965347997168294   0.3907536210162571   0.19332053721474513   0.24935243703686755   0.8494941990738512   0.6341589075279351   0.33840762339308883   0.4586354510850482   0.21496237167385124   0.6150137486113473   0.9396727205696299   0.7292323498454217   0.11906337489496852   0.8792163596930791   0.46029151986473116   0.3202236876590435   0.12645137797274333   0.7985373211178851   0.14153055065323888   0.06527597559657465   0.031604609949409626   0.7332868154879078   0.054768901746892196   0.9465948898122405   0.1350698102325803   0.34253319447165065   0.861448364532147   0.6972424527753729   0.2855756111587291   0.7083742869437155   0.5230407411390582   0.23860700169032473   0.07061323948487788   0.09336053833236822   0.5833680205694284   0.5093746518449029   0.9515498645899093   0.21414417863928914   0.12307650070469717   0.18915096418585944   0.825098486617166   0.415606857521404   0.9815459500514583   0.12387498858928478   0.7934938766677564
0.6823200420334963   0.9267770483045661   0.17728009877704431   0.6584240664351761   0.33978684756184563   0.06532868377241904   0.48003764600167137   0.372848455276447   0.6314125606181301   0.5422879426333608   0.24143064431134667   0.3022352157915691   0.5380520222857619   0.9589199220639325   0.7320559924664437   0.3506853512016598   0.32390784364647274   0.8358434213592353   0.5429050282805843   0.5255868645844938   0.9083009861250687   0.854297471307777   0.4190300396912995   0.7320929879167374   0.22598094409157246   0.9275204230032109   0.24174994091425517   0.07366892148156122   0.8861940965297268   0.862191739230792   0.7617122949125839   0.7008204662051143   0.25478153591159675   0.31990379659743107   0.5202816506012371   0.39858525041354514   0.7167295136258348   0.36098387453349856   0.7882256581347934   0.04789989921188537   0.3928216699793621   0.5251404531742633   0.2453206298542092   0.5223130346273916   0.48452068385429337   0.6708429818664862   0.8262905901629097   0.7902200467106543   0.2585397397627209   0.7433225588632753   0.5845406492486546   0.7165511252290931   0.372345643232994   0.8811308196324834   0.8228283543360707   0.015730659023978855   0.1175641073213973   0.5612270230350523   0.3025467037348336   0.6171454086104338   0.40083459369556246   0.20024314850155372   0.5143210456000401   0.5692455093985483
0.008012923716200404   0.6751026953272905   0.26900041574583095   0.04693247477115672   0.5234922398619071   0.004259713460804254   0.44270982558292127   0.2567124280605024   0.2649525000991862   0.260937154597529   0.8581691763342667   0.5401613028314093   0.8926068568661921   0.3798063349650456   0.03534082199819599   0.5244306438074304   0.7750427495447949   0.8185793119299933   0.7327941182633624   0.9072852351969968   0.3742081558492324   0.6183361634284396   0.21847307266332225   0.3380397257984484   0.36619523213303196   0.943233468101149   0.9494726569174913   0.2911072510272916   0.8427029922711249   0.9389737546403448   0.50676283133457   0.034394822966789244   0.5777504921719387   0.6780366000428159   0.6485936550003033   0.4942335201353799   0.6851436353057466   0.2982302650777703   0.6132528330021073   0.9698028763279495   0.9101008857609517   0.47965095314777695   0.8804587147387449   0.06251764113095276   0.5358927299117193   0.8613147897193374   0.6619856420754227   0.7244779153325044   0.16969749777868737   0.9180813216181882   0.7125129851579314   0.43337066430521276   0.3269945055075624   0.9791075669778434   0.20575015382336131   0.3989758413384235   0.7492440133356237   0.30107096693502755   0.557156498823058   0.9047423212030435   0.06410037802987711   0.002840701857257292   0.9439036658209506   0.9349394448750941
0.15399949226892537   0.5231897487094803   0.06344495108220573   0.8724218037441414   0.6181067623572061   0.6618749589901429   0.40145930900678306   0.14794388841163694   0.44840926457851865   0.7437936373719547   0.6889463238488517   0.7145732241064242   0.12141475907095624   0.7646860703941112   0.48319617002549037   0.31559738276800064   0.37217074573533254   0.4636151034590837   0.9260396712024324   0.4108550615649571   0.30807036770545543   0.46077440160182637   0.9821360053814817   0.475915616689863   0.15407087543653006   0.937584652892346   0.918691054299276   0.6034938129457217   0.535964113079324   0.2757096939022031   0.5172317452924929   0.4555499245340847   0.08755484850080533   0.5319160565302484   0.8282854214436413   0.7409767004276605   0.9661400894298491   0.7672299861361372   0.3450892514181509   0.42537931765965986   0.5939693436945166   0.30361488267705355   0.41904958021571853   0.014524256094702783   0.2858989759890611   0.8428404810752272   0.4369135748342368   0.5386086394048398   0.13182810055253108   0.9052558281828812   0.5182225205349609   0.9351148264591181   0.5958639874732071   0.6295461342806781   0.0009907752424679567   0.47956490192503337   0.5083091389724017   0.09763007775042959   0.17270535379882673   0.7385882014973728   0.5421690495425526   0.33040009161429235   0.8276161023806758   0.31320888383771295
0.9481997058480361   0.026785208937238788   0.4085665221649573   0.29868462774301013   0.6623007298589749   0.1839447278620116   0.9716529473307205   0.7600759883381704   0.5304726293064439   0.27868889967913046   0.4534304267957596   0.8249611618790522   0.9346086418332368   0.6491427653984524   0.4524396515532917   0.3453962599540189   0.426299502860835   0.5515126876480229   0.27973429775446496   0.6068080584566461   0.8841304533182823   0.22111259603373046   0.4521181953737891   0.29359917461893315   0.9359307474702463   0.1943273870964917   0.04355167320883176   0.994914546875923   0.2736300176112713   0.010382659234480089   0.07189872587811125   0.2348385585377526   0.7431573883048275   0.7316937595553497   0.6184682990823516   0.4098773966587003   0.8085487464715907   0.08255099415689723   0.1660286475290599   0.06448113670468143   0.38224924361075563   0.5310383065088744   0.886294349774595   0.4576730782480354   0.49811879029247325   0.30992571047514395   0.43417615440080587   0.16407390362910224   0.562188042822227   0.11559832337865225   0.39062448119197407   0.16915935675317925   0.28855802521095564   0.10521566414417216   0.3187257553138628   0.9343207982154267   0.5454006369061282   0.3735219045888225   0.7002574562315113   0.5244434015567263   0.7368518904345375   0.2909709104319253   0.5342288087024513   0.4599622648520449
0.35460264682378184   0.7599326039230508   0.6479344589278564   0.0022891866040095276   0.8564838565313087   0.45000689344790695   0.21375830452705052   0.8382152829749073   0.29429581370908164   0.3344085700692547   0.8231338233350765   0.669055926221728   0.005737788498125993   0.22919290592508254   0.5044080680212136   0.7347351280063014   0.4603371515919978   0.8556710013362601   0.8041506117897024   0.21029172644957503   0.7234852611574603   0.5647000909043347   0.2699218030872511   0.7503294615975301   0.3688826143336784   0.8047674869812839   0.6219873441593947   0.7480402749935205   0.5123987578023699   0.3547605935333769   0.4082290396323442   0.9098249920186133   0.2181029440932882   0.020352023464122192   0.5850952162972678   0.24076906579688528   0.2123651555951622   0.7911591175390397   0.08068714827605417   0.5060339377905839   0.7520280040031644   0.9354881162027796   0.2765365364863518   0.2957422113410089   0.028542742845704086   0.3707880252984449   0.006614733399100684   0.5454127497434788   0.6596601285120256   0.566020538317161   0.38462738923970596   0.7973724747499582   0.1472613707096558   0.21125994478378418   0.9763983496073617   0.8875474827313449   0.9291584266163676   0.19090792131966197   0.391303133310094   0.6467784169344596   0.7167932710212054   0.39974880378062233   0.3106159850340398   0.14074447914387567
0.964765267018041   0.46426068757784267   0.03407944854768802   0.8450022678028668   0.936222524172337   0.09347266227939778   0.027464715148587334   0.299589518059388   0.2765623956603113   0.5274521239622367   0.6428373259088814   0.5022170433094298   0.12930102495065549   0.31619217917845255   0.6664389763015196   0.6146695605780849   0.20014259833428785   0.12528425785879055   0.2751358429914257   0.9678911436436253   0.48334932731308244   0.7255354540781682   0.9645198579573859   0.8271466644997496   0.5185840602950414   0.26127476650032555   0.9304404094096979   0.9821443966968828   0.5823615361227045   0.16780210422092776   0.9029756942611106   0.6825548786374949   0.30579914046239315   0.640349980258691   0.26013836835222914   0.18033783532806508   0.1764981155117377   0.3241578010802385   0.5936993920507095   0.5656682747499802   0.9763555171774498   0.19887354322144793   0.31856354905928386   0.5977771311063549   0.4930061898643674   0.4733380891432797   0.35404369110189793   0.7706304666066053   0.974422129569326   0.21206332264295416   0.4236032816922001   0.7884860699097224   0.3920605934466215   0.04426121842202641   0.5206275874310895   0.10593119127222753   0.08626145298422833   0.40391123816333535   0.26048921907886036   0.9255933559441625   0.9097633374724906   0.07975343708309689   0.6667898270281508   0.3599250811941823
0.9334078202950408   0.880879893861649   0.34822627796886696   0.7621479500878274   0.44040163043067343   0.40754180471836926   0.994182586866969   0.9915174834812222   0.4659795008613475   0.1954784820754151   0.570579305174769   0.2030314135714998   0.07391890741472597   0.1512172636533887   0.04995171774367948   0.09710022229927229   0.9876574544304977   0.7473060254900533   0.7894624986648191   0.17150686635510984   0.07789411695800699   0.6675525884069564   0.12267267163666834   0.8115817851609275   0.14448629666296617   0.7866726945453074   0.7744463936678013   0.04943383507310011   0.7040846662322927   0.3791308898269382   0.7802638068008323   0.05791635159187792   0.23810516537094528   0.1836524077515231   0.20968450162606334   0.8548849380203781   0.16418625795621933   0.03243514409813442   0.15973278388238385   0.7577847157211058   0.1765288035257217   0.2851291186080811   0.3702702852175647   0.586277849365996   0.0986346865677147   0.6175765302011247   0.24759761358089638   0.7746960642050684   0.9541483899047485   0.8309038356558173   0.473151219913095   0.7252622291319684   0.2500637236724558   0.45177294582887906   0.6928874131122627   0.6673458775400904   0.011958558301510474   0.2681205380773559   0.48320291148619937   0.8124609395197123   0.8477723003452912   0.2356853939792215   0.3234701276038155   0.054676223798606476
0.6712434968195695   0.9505562753711404   0.9531998423862508   0.46839837443261045   0.5726088102518547   0.3329797451700157   0.7056022288053544   0.693702310227542   0.6184604203471062   0.5020759095141984   0.23245100889225936   0.9684400810955737   0.3683966966746505   0.05030296368531943   0.5395635957799967   0.3010942035554833   0.35643813837314003   0.7821824256079635   0.05636068429379732   0.48863326403577095   0.5086658380278489   0.546497031628742   0.7328905566899818   0.43395704023716447   0.8374223412082794   0.5959407562576016   0.779690714303731   0.965558665804554   0.2648135309564246   0.2629610110875859   0.07408848549837667   0.271856355577012   0.6463531106093183   0.7608851015733874   0.8416374766061173   0.3034162744814383   0.27795641393466786   0.710582137888068   0.30207388082612063   0.0023220709259550425   0.9215182755615279   0.9283997122801045   0.2457131965323233   0.513688806890184   0.41285243753367895   0.3819026806513625   0.5128226398423414   0.0797317666530196   0.5754300963253995   0.7859619243937609   0.7331319255386104   0.1141731008484656   0.3106165653689749   0.523000913306175   0.6590434400402337   0.8423167452714536   0.6642634547596565   0.7621158117327876   0.8174059634341164   0.5389004707900154   0.3863070408249887   0.0515336738447196   0.5153320826079958   0.5365783998640603
0.4647887652634608   0.1231339615646151   0.2696188860756725   0.022889592973876192   0.05193632772978184   0.7412312809132526   0.7567962462333311   0.9431578263208565   0.47650623140438225   0.9552693565194917   0.023664320694720638   0.828984725472391   0.16588966603540733   0.43226844321331664   0.3646208806544869   0.9866679802009374   0.5016262112757508   0.6701526314805291   0.5472149172203704   0.447767509410922   0.11531917045076213   0.6186189576358094   0.03188283461237465   0.9111891095468617   0.6505304051873013   0.49548499607119434   0.7622639485367021   0.8882995165729856   0.5985940774575195   0.7542537151579417   0.00546770230337109   0.945141690252129   0.12208784605313722   0.7989843586384501   0.9818033816086504   0.116156964779738   0.9561981800177298   0.3667159154251334   0.6171825009541636   0.12948898457880065   0.4545719687419791   0.6965632839446043   0.06996758373379308   0.6817214751678786   0.33925279829121696   0.07794432630879487   0.03808474912141844   0.7705323656210169   0.6887223931039156   0.5824593302376005   0.2758208005847163   0.8822328490480313   0.09012831564639612   0.8282056150796587   0.27035309828134524   0.9370911587959023   0.9680404695932588   0.029221256441208713   0.28854971667269474   0.8209341940161643   0.011842289575529017   0.6625053410160753   0.6713672157185312   0.6914452094373637
0.55727032083355   0.965942057071471   0.6013996319847381   0.00972373426948505   0.218017522542333   0.8879977307626761   0.5633148828633197   0.23919136864846818   0.5292951294384174   0.3055384005250756   0.2874940822786034   0.3569585196004369   0.43916681379202127   0.47733278544541685   0.017140983997258167   0.4198673608045346   0.47112634419876237   0.44811152900420814   0.7285912673245634   0.5989331667883703   0.45928405462323335   0.7856061879881328   0.057224051606032195   0.9074879573510065   0.9020137337896834   0.8196641309166618   0.45582441962129405   0.8977642230815215   0.6839962112473504   0.9316664001539857   0.8925095367579744   0.6585728544330534   0.15470108180893302   0.6261279996289101   0.605015454479371   0.30161433483261646   0.7155342680169118   0.14879521418349326   0.5878744704821128   0.8817469740280819   0.24440792381814935   0.7006836851792851   0.8592832031575495   0.28281380723971167   0.785123869194916   0.9150774971911524   0.8020591515515172   0.3753258498887051   0.8831101354052325   0.09541336627449053   0.3462347319302232   0.4775616268071836   0.19911392415788212   0.16374696612050482   0.4537251951722488   0.8189887723741303   0.044412842348949114   0.5376189664915947   0.8487097406928777   0.5173744375415138   0.3288785743320374   0.38882375230810146   0.2608352702107649   0.6356274635134319
0.08447065051388802   0.6881400671288164   0.4015520670532155   0.35281365627372024   0.2993467813189721   0.773062569937664   0.5994929155016983   0.9774878063850152   0.4162366459137395   0.6776492036631735   0.25325818357147506   0.4999261795778316   0.21712272175585737   0.5139022375426686   0.7995329883992263   0.6809374072037013   0.17270987940690824   0.9762832710510739   0.9508232477063485   0.16356296966218747   0.8438313050748709   0.5874595187429724   0.6899879774955836   0.5279355061487556   0.7593606545609828   0.899319451614156   0.2884359104423681   0.1751218498750353   0.46001387324201076   0.12625688167649207   0.6889429949406699   0.19763404349002014   0.043777227328271294   0.4486076780133186   0.4356848113691948   0.6977078639121885   0.8266545055724139   0.93470544047065   0.6361518229699685   0.01677045670848727   0.6539446261655056   0.958422169419576   0.68532857526362   0.8532074870462998   0.8101133210906348   0.3709626506766036   0.9953405977680364   0.3252719808975442   0.050752666529651984   0.47164319906244756   0.7069046873256682   0.15015013102250893   0.5907387932876412   0.34538631738595543   0.017961692384998427   0.9525160875324887   0.54696156595937   0.8967786393726368   0.5822768810158037   0.2548082236203002   0.720307060386956   0.9620731989019868   0.9461250580458351   0.23803776691181294
0.06636243422145029   0.003651029482410838   0.2607964827822151   0.38483027986551316   0.25624911313081544   0.6326883788058072   0.2654558850141787   0.05955829896796893   0.20549644660116348   0.1610451797433597   0.5585511976885105   0.90940816794546   0.6147576533135223   0.8156588623574043   0.540589505303512   0.9568920804129712   0.06779608735415239   0.9188802229847673   0.9583126242877084   0.702083856792671   0.3474890269671964   0.9568070240827805   0.01218756624187325   0.4640460898808581   0.28112659274574614   0.9531559946003697   0.7513910834596581   0.07921581001534495   0.02487747961493066   0.32046761579456245   0.4859351984454794   0.01965751104737601   0.8193810330137672   0.15942243605120276   0.927384000756969   0.11024934310191599   0.20462337970024488   0.3437635736937985   0.38679449545345695   0.15335726268894476   0.13682729234609248   0.42488335070903116   0.4284818711657486   0.45127340589627374   0.7893382653788961   0.46807632662625065   0.41629430492387537   0.9872273160154157   0.5082116726331499   0.514920332025881   0.6649032214642172   0.9080115060000707   0.4833341930182193   0.19445271623131852   0.17896802301873782   0.8883539949526947   0.6639531600044521   0.03503028018011575   0.25158402226176885   0.7781046518507787   0.45932978030420724   0.6912667064863173   0.8647895268083119   0.6247473891618339
0.32250248795811476   0.26638335577728606   0.43630765564256324   0.1734739832655602   0.5331642225792187   0.7983070291510355   0.020013350718687907   0.18624666725014458   0.024952549946068738   0.28338669712515446   0.35511012925447066   0.27823516125007386   0.5416183569278494   0.08893398089383596   0.17614210623573284   0.3898811662973792   0.8776651969233974   0.05390370071372021   0.924558083973964   0.6117765144466005   0.4183354166191901   0.362636994227403   0.05976855716565211   0.9870291252847666   0.09583292866107537   0.0962536384501169   0.6234609015230889   0.8135551420192063   0.5626687060818567   0.29794660929908146   0.6034475508044009   0.6273084747690618   0.5377161561357879   0.014559912173926983   0.24833742154993027   0.3490733135189879   0.9960977992079385   0.9256259312800911   0.07219531531419743   0.9591921472216087   0.11843260228454115   0.8717222305663708   0.14763723134023343   0.3474156327750082   0.7000971856653511   0.5090852363389679   0.08786867417458133   0.36038650749024165   0.6042642570042757   0.41283159788885093   0.46440777265149247   0.5468313654710353   0.04159555092241897   0.11488498858976946   0.8609602218470915   0.9195228907019736   0.503879394786631   0.10032507641584247   0.6126228002971613   0.5704495771829856   0.5077815955786925   0.17469914513575147   0.5404274849829639   0.6112574299613769
0.38934899329415135   0.30297691456938064   0.3927902536427304   0.26384179718636874   0.6892518076288003   0.7938916782304128   0.3049215794681491   0.9034552896961271   0.08498755062452466   0.38106008034156186   0.8405138068166566   0.35662392422509176   0.0433919997021057   0.26617509175179244   0.979553584969565   0.43710103352311824   0.5395126049154747   0.16585001533594995   0.36693078467240375   0.8666514563401326   0.031731009336782176   0.9911508702001985   0.8265032996894399   0.2553940263787557   0.6423820160426308   0.6881739556308178   0.4337130460467095   0.991552229192387   0.9531302084138304   0.894282277400405   0.12879146657856042   0.0880969394962599   0.8681426577893059   0.5132221970588432   0.28827765976190384   0.7314730152711681   0.8247506580872002   0.24704710530705074   0.30872407479233877   0.2943719817480499   0.28523805317172546   0.0811970899711008   0.941793290119935   0.4277205254079173   0.25350704383494327   0.09004621977090231   0.11528999043049507   0.1723264990291616   0.6111250277923125   0.4018722641400844   0.6815769443837856   0.18077426983677466   0.6579948193784819   0.5075899867396794   0.5527854778052251   0.09267733034051477   0.7898521615891761   0.9943677896808363   0.2645078180433213   0.36120431506934664   0.965101503501976   0.7473206843737855   0.9557837432509826   0.06683233332129675
0.6798634503302505   0.6661235944026846   0.013990453131047558   0.6391118079133794   0.42635640649530726   0.5760773746317823   0.8987004627005525   0.4667853088842178   0.8152313787029948   0.17420511049169793   0.21712351831676693   0.2860110390474432   0.1572365593245129   0.6666151237520185   0.6643380405115418   0.1933337087069284   0.36738439773533677   0.6722473340711823   0.3998302224682205   0.8321293936375818   0.4022828942333608   0.9249266496973968   0.4440464792172379   0.765297060316285   0.7224194439031102   0.25880305529471215   0.43005602608619037   0.12618525240290554   0.29606303740780293   0.6827256806629298   0.5313555633856378   0.6593999435186877   0.48083165870480815   0.5085205701712319   0.3142320450688709   0.37338890447124456   0.32359509938029524   0.8419054464192133   0.6498940045573292   0.18005519576431614   0.9562107016449585   0.16965811234803102   0.2500637820891087   0.3479258021267344   0.5539278074115978   0.24473146265063422   0.8060173028718708   0.5826287418104494   0.8315083635084874   0.985928407355922   0.3759612767856804   0.45644348940754387   0.5354453261006845   0.3032027266929923   0.8446057134000425   0.7970435458888562   0.054613667395876406   0.7946821565217604   0.5303736683311716   0.42365464141761155   0.7310185680155812   0.9527767101025472   0.8804796637738425   0.24359944565329542
0.7748078663706226   0.7831185977545161   0.6304158816847337   0.895673643526561   0.22088005895902493   0.5383871351038819   0.8243985788128629   0.31304490171611166   0.3893716954505374   0.5524587277479598   0.4484373020271825   0.8566014123085678   0.8539263693498529   0.2492560010549675   0.6038315886271399   0.05955786641971167   0.7993127019539765   0.45457384453320704   0.07345792029596832   0.6359032250021001   0.06829413393839531   0.50179713443066   0.19297825652212583   0.39230377934880467   0.2934862675677727   0.7186785366761438   0.562562374837392   0.49663013582224363   0.07260620860874775   0.18029140157226195   0.7381637960245291   0.183585234106132   0.6832345131582104   0.6278326738243021   0.2897264939973465   0.32698382179756424   0.8293081438083575   0.3785766727693346   0.6858949053702066   0.2674259553778526   0.029995441854380977   0.9240028282361276   0.6124369850742383   0.6315227303757525   0.9617013079159856   0.42220569380546763   0.4194587285521124   0.2392189510269478   0.668215040348213   0.7035271571293238   0.8568963537147204   0.7425888152047041   0.5956088317394652   0.5232357555570618   0.11873255769019128   0.5590035810985721   0.912374318581255   0.8954030817327597   0.8290060636928448   0.23201975930100788   0.08306617477289746   0.5168264089634251   0.14311115832263818   0.9645938039231553
0.05307073291851648   0.5928235807272976   0.5306741732483999   0.3330710735474029   0.09136942500253083   0.17061788692182994   0.11121544469628754   0.0938521225204551   0.4231543846543178   0.46709072979250615   0.2543190909815672   0.351263307315751   0.8275455529148525   0.9438549742354443   0.13558653329137588   0.7922597262171789   0.9151712343335977   0.0484518925026846   0.30658046959853114   0.560239966916171   0.8321050595607002   0.5316254835392595   0.16346931127589293   0.5956461629930156   0.7790343266421837   0.938801902811962   0.632795138027493   0.26257508944561275   0.6876649016396529   0.7681840158901321   0.5215796933312055   0.16872296692515765   0.26451051698533506   0.30109328609762587   0.2672606023496383   0.8174596596094067   0.43696496407048246   0.3572383118621816   0.1316740690582624   0.025199933392227782   0.5217937297368848   0.30878641935949697   0.8250935994597313   0.4649599664760568   0.6896886701761845   0.7771609358202375   0.6616242881838383   0.8693138034830412   0.9106543435340008   0.8383590330082755   0.02882915015634533   0.6067387140374284   0.2229894418943479   0.0701750171181435   0.5072494568251399   0.43801574711227076   0.9584789249090129   0.7690817310205176   0.23998885447550158   0.6205560875028642   0.5215139608385303   0.41184341915833605   0.1083147854172392   0.5953561541106364
0.9997202311016455   0.10305699979883907   0.28322118595750795   0.13039618763457952   0.31003156092546097   0.3258960639786016   0.6215968977736697   0.2610823841515384   0.39937721739146015   0.4875370309703261   0.5927677476173243   0.65434367011411   0.17638777549711226   0.4173620138521826   0.08551829079218441   0.21632792300183917   0.21790885058809945   0.648280282831665   0.8455294363166829   0.595771835498975   0.6963948897495691   0.2364368636733289   0.7372146508994436   0.00041568138833872445   0.6966746586479236   0.1333798638744898   0.45399346494193565   0.8700194937537592   0.3866430977224626   0.8074837998958883   0.832396567168266   0.6089371096022208   0.9872658803310024   0.3199467689255621   0.23962881955094176   0.9545934394881108   0.8108781048338901   0.9025847550733795   0.15411052875875733   0.7382655164862717   0.5929692542457907   0.25430447224171465   0.30858109244207454   0.14249368098729662   0.8965743644962215   0.017867608568385738   0.5713664415426309   0.1420779995989579   0.199899705848298   0.8844877446938959   0.11737297660069523   0.2720585058451987   0.8132566081258354   0.07700394479800772   0.2849764094324292   0.6631213962429778   0.8259907277948331   0.7570571758724456   0.04534758988148742   0.708527956754867   0.015112622960942922   0.854472420799066   0.89123706112273   0.9702624402685953
0.42214336871515223   0.6001679485573514   0.5826559686806556   0.8277687592812987   0.5255690042189307   0.5823003399889657   0.011289527138024657   0.6856907596823408   0.3256692983706327   0.6978125952950698   0.8939165505373294   0.41363225383714214   0.5124126902447972   0.620808650497062   0.6089401411049002   0.7505108575941642   0.6864219624499642   0.8637514746246164   0.5635925512234128   0.041982900839297226   0.6713093394890213   0.0092790538255504   0.6723554901006827   0.07172046057070189   0.249165970773869   0.409111105268199   0.08969952142002718   0.24395170128940316   0.7235969665549383   0.8268107652792334   0.07840999428200253   0.5582609416070623   0.39792766818430564   0.1289981699841636   0.1844934437446731   0.1446286877699202   0.8855149779395084   0.5081895194871016   0.5755533026397729   0.39411783017575597   0.19909301548954425   0.6444380448624852   0.011960751416360032   0.35213492933645874   0.527783676000523   0.6351589910369347   0.3396052613156773   0.2804144687657568   0.27861770522665397   0.2260478857687358   0.2499057398956501   0.03646276747635368   0.5550207386717156   0.39923712048950244   0.17149574561364758   0.47820182586929133   0.15709307048740997   0.2702389505053388   0.9870023018689744   0.33357313809937117   0.27157809254790155   0.7620494310182372   0.4114489992292016   0.9394553079236152
0.0724850770583573   0.11761138615575202   0.3994882478128416   0.5873203785871565   0.5447014010578343   0.4824523951188172   0.05988298649716429   0.30690590982139965   0.2660836958311803   0.2564045093500814   0.8099772466015142   0.27044314234504596   0.7110629571594647   0.857167388860579   0.6384815009878666   0.7922413164757547   0.5539698866720547   0.5869284383552401   0.6514791991188922   0.45866817837638346   0.28239179412415316   0.8248790073370029   0.24003019988969054   0.5192128704527682   0.20990671706579583   0.707267621181251   0.840541952076849   0.9318924918656117   0.6652053160079615   0.2248152260624337   0.7806589655796847   0.6249865820442121   0.3991216201767812   0.9684107167123522   0.9706817189781705   0.35454343969916613   0.6880586630173166   0.1112433278517733   0.33220021799030386   0.5623021232234114   0.13408877634526187   0.5243148894965332   0.6807210188714117   0.103633944847028   0.8516969822211087   0.6994358821595301   0.4406908189817212   0.5844210743942597   0.6417902651553129   0.9921682609782793   0.6001488669048722   0.652528582528648   0.9765849491473514   0.7673530349158455   0.8194899013251875   0.027542000484435877   0.5774633289705701   0.7989423182034933   0.848808182347017   0.6729985607852698   0.8894046659532535   0.68769899035172   0.5166079643567132   0.11069643756185829
0.7553158896079917   0.16338410085518681   0.8358869454853014   0.007062492714830297   0.903618907386883   0.46394821869565667   0.39519612650358027   0.42264141832057056   0.2618286422315701   0.4717799577173774   0.795047259598708   0.7701128357919226   0.28524369308421876   0.704426922801532   0.9755573582735205   0.7425708353074867   0.7077803641136486   0.9054846045980387   0.12674917592650353   0.06957227452221694   0.8183756981603951   0.21778561424631873   0.6101412115697904   0.9588758369603586   0.0630598085524034   0.05440151339113191   0.7742542660844889   0.9518133442455283   0.1594409011655204   0.5904532946954753   0.37905813958090867   0.5291719259249578   0.8976122589339504   0.11867333697809783   0.5840108799822006   0.7590590901330352   0.6123685658497315   0.4142464141765659   0.6084535217086801   0.0164882548255485   0.9045882017360829   0.5087618095785272   0.4817043457821765   0.9469159803033316   0.08621250357568778   0.2909761953322085   0.8715631342123862   0.988040143342973   0.0231526950232844   0.2365746819410766   0.09730886812789721   0.036226799097444584   0.863711793857764   0.6461213872456013   0.7182507285469886   0.5070548731724868   0.9660995349238137   0.5274480502675035   0.134239848564788   0.7479957830394516   0.35373096907408214   0.11320163609093759   0.5257863268561079   0.7315075282139031
0.4491427673379993   0.6044398265124103   0.044081981073931464   0.7845915479105715   0.36293026376231147   0.3134636311802019   0.17251884686154534   0.7965514045675987   0.3397775687390271   0.0768889492391253   0.07520997873364813   0.760324605470154   0.47606577488126306   0.430767561993524   0.3569592501866596   0.2532697322976672   0.5099662399574494   0.9033195117260205   0.22271940162187157   0.5052739492582157   0.15623527088336725   0.790117875635083   0.6969330747657636   0.7737664210443125   0.707092503545368   0.18567804912267255   0.6528510936918321   0.989174873133741   0.3441622397830565   0.8722144179424707   0.4803322468302868   0.19262346856614238   0.004384671044029433   0.7953254687033453   0.4051222680966387   0.43229886309598836   0.5283188961627664   0.36455790670982136   0.04816301790997913   0.1790291307983211   0.01835265620531695   0.46123839498380087   0.8254436162881076   0.6737551815401055   0.8621173853219497   0.671120519348718   0.12851054152234395   0.899988760495793   0.15502488177658172   0.4854424702260454   0.47565944783051184   0.910813887362052   0.8108626419935252   0.6132280522835748   0.995327201000225   0.7181904187959096   0.8064779709494958   0.8179025835802294   0.5902049329035863   0.2858915556999213   0.2781590747867294   0.4533446768704081   0.5420419149936072   0.10686242490160017
0.25980641858141246   0.9921062818866072   0.7165982987054996   0.43310724336149464   0.39768903325946275   0.32098576253788924   0.5880877571831556   0.5331184828657016   0.24266415148288106   0.8355432923118438   0.11242830935264386   0.6223045955036497   0.43180150948935586   0.22231524002826902   0.11710110835241885   0.9041141767077401   0.6253235385398601   0.4044126564480396   0.5268961754488325   0.6182226210078188   0.34716446375313065   0.9510679795776316   0.9848542604552253   0.5113601961062185   0.08735804517171818   0.9589616976910244   0.26825596174972566   0.0782529527447239   0.6896690119122554   0.6379759351531351   0.68016820456657   0.5451344698790223   0.4470048604293744   0.8024326428412913   0.5677398952139261   0.9228298743753726   0.015203350940018494   0.5801174028130224   0.45063878686150727   0.01871569766763251   0.3898798124001584   0.17570474636498273   0.9237426114126748   0.40049307665981376   0.04271534864702776   0.22463676678735117   0.9388883509574495   0.8891328805535952   0.9553573034753096   0.2656750690963268   0.6706323892077238   0.8108799278088713   0.2656882915630542   0.6276991339431917   0.9904641846411538   0.2657454579298491   0.8186834311336798   0.8252664911019003   0.4227242894272277   0.3429155835544766   0.8034800801936614   0.24514908828887802   0.9720855025657203   0.32419988588684406
0.4136002677935029   0.06944434192389529   0.04834289115304563   0.9237068092270303   0.37088491914647514   0.8448075751365441   0.10945454019559618   0.03457392867343507   0.4155276156711656   0.5791325060402173   0.4388221509878724   0.22369400086456373   0.1498393241081114   0.9514333720970256   0.4483579663467186   0.9579485429347147   0.3311558929744316   0.12616688099512527   0.025633676919490943   0.615032959380238   0.5276758127807702   0.8810177927062472   0.05354817435377055   0.290833073493394   0.11407554498726737   0.811573450782352   0.005205283200724917   0.3671262642663637   0.7431906258407922   0.9667658756458078   0.8957507430051287   0.3325523355929286   0.3276630101696266   0.3876333696055906   0.45692859201725633   0.10885833472836487   0.17782368606151522   0.436199997508565   0.008570625670537714   0.15090979179365024   0.8466677930870836   0.3100331165134397   0.9829369487510468   0.5358768324134122   0.31899198030631337   0.42901532380719243   0.9293887743972762   0.24504375892001826   0.204916435319046   0.6174418730248404   0.9241834911965513   0.8779174946536545   0.46172580947825376   0.6506759973790326   0.02843274819142257   0.545365159060726   0.13406279930862713   0.26304262777344195   0.5715041561741663   0.4365068243323611   0.956239113247112   0.826842630264877   0.5629335305036285   0.2855970325387109
0.1095713201600283   0.5168095137514374   0.5799965817525817   0.7497202001252986   0.790579339853715   0.08779418994424491   0.6506078073553055   0.5046764412052804   0.585662904534669   0.4703523169194045   0.7264243161587542   0.6267589465516258   0.1239370950564152   0.8196763195403719   0.6979915679673316   0.08139378749089986   0.9898742957477881   0.55663369176693   0.12648741179316542   0.6448869631585388   0.033635182500676146   0.729791061502053   0.5635538812895369   0.3592899306198279   0.9240638623406479   0.21298154775061565   0.9835572995369551   0.6095697304945292   0.1334845224869329   0.12518735780637075   0.3329494921816496   0.10489328928924885   0.5478216179522639   0.6548350408869663   0.6065251760228954   0.478134342737623   0.4238845228958487   0.8351587213465943   0.9085336080555637   0.39674055524672314   0.43401022714806065   0.27852502957966435   0.7820461962623982   0.7518535920881844   0.4003750446473845   0.5487339680776114   0.21849231497286137   0.39256366146835653   0.47631118230673664   0.3357524203269957   0.23493501543590622   0.7829939309738273   0.34282665981980376   0.21056506252062498   0.9019855232542566   0.6781006416845784   0.7950050418675398   0.5557300216336587   0.2954603472313613   0.19996629894695542   0.3711205189716911   0.7205713002870644   0.38692673917579756   0.8032257437002323
0.9371102918236305   0.44204627070740005   0.6048805429133993   0.05137215161204784   0.536735247176246   0.8933123026297887   0.38638822794053795   0.6588084901436914   0.06042406486950934   0.557559882302793   0.1514532125046317   0.8758145591698641   0.7175974050497056   0.34699481978216795   0.24946768925037507   0.19771391748528563   0.9225923631821658   0.7912647981485093   0.9540073420190138   0.9977476185383302   0.5514718442104746   0.07069349786144485   0.5670806028432163   0.19452187483809796   0.6143615523868441   0.6286472271540449   0.9622000599298169   0.14314972322605013   0.07762630521059814   0.7353349245242562   0.575811831989279   0.48434123308235877   0.017202240341088804   0.17777504222146326   0.42435861948464726   0.6085266739124947   0.2996048352913832   0.8307802224392953   0.1748909302342722   0.4108127564272091   0.37701247210921746   0.03951542429078608   0.2208835882152584   0.41306513788887894   0.8255406278987428   0.9688219264293412   0.6538029853720422   0.21854326305078095   0.2111790755118987   0.3401746992752964   0.6916029254422252   0.07539353982473083   0.13355277030130058   0.6048397747510402   0.11579109345294623   0.5910523067423721   0.11635052996021178   0.42706473252957694   0.691432473968299   0.9825256328298773   0.8167456946688285   0.5962845100902816   0.5165415437340267   0.5717128764026682
0.43973322255961106   0.5567690857994956   0.2956579555187684   0.15864773851378924   0.6141925946608682   0.5879471593701543   0.6418549701467262   0.9401044754630083   0.4030135191489695   0.2477724600948579   0.950252044704501   0.8647109356382775   0.2694607488476689   0.6429326853438178   0.8344609512515547   0.2736586288959054   0.15311021888745716   0.21586795281424076   0.1430284772832558   0.2911329960660281   0.3363645242186286   0.6195834427239592   0.626486933549229   0.71942011966336   0.8966313016590175   0.06281435692446362   0.3308289780304607   0.5607723811495707   0.28243870699814927   0.4748671975543093   0.6889740078837344   0.6206679056865624   0.8794251878491798   0.22709473745945138   0.7387219631792334   0.7559569700482849   0.6099644390015109   0.5841620521156337   0.9042610119276787   0.4822983411523795   0.4568542201140537   0.36829409930139295   0.761232534644423   0.19116534508635138   0.1204896958954251   0.7487106565774337   0.1347456010951939   0.4717452254229914   0.22385839423640758   0.6858962996529702   0.8039166230647332   0.9109728442734207   0.9414196872382583   0.21102910209866085   0.11494261518099876   0.29030493858685835   0.061994499389078514   0.9839343646392095   0.3762206520017653   0.5343479685385734   0.45203006038756766   0.39977231252357576   0.47195964007408653   0.05204962738619389
0.9951758402735139   0.031478213222182846   0.7107271054296636   0.8608842822998425   0.8746861443780889   0.28276755664474906   0.5759815043344697   0.3891390568768511   0.6508277501416813   0.5968712569917789   0.7720648812697365   0.47816621260343034   0.709408062903423   0.385842154893118   0.6571222660887377   0.187861274016572   0.6474135635143444   0.40190779025390855   0.2809016140869724   0.6535133054779986   0.1953835031267768   0.0021354777303327953   0.8089419740128859   0.6014636780918047   0.20020766285326283   0.9706572645081499   0.0982148685832223   0.7405793957919622   0.32552151847517397   0.6878897078634009   0.5222333642487527   0.3514403389151111   0.6746937683334927   0.091018450871622   0.7501684829790162   0.8732741263116808   0.9652857054300698   0.705176295978504   0.09304621689027846   0.6854128522951088   0.31787214191572527   0.3032685057245954   0.812144602803306   0.031899546817110214   0.12248863878894847   0.3011330279942626   0.0032026287904201576   0.4304358687253055   0.9222809759356856   0.33047576348611263   0.9049877602071978   0.6898564729333433   0.5967594574605116   0.6425860556227118   0.38275439595844524   0.3384161340182322   0.9220656891270189   0.5515676047510898   0.6325859129794291   0.46514200770655134   0.9567799836969492   0.8463913087725858   0.5395396960891506   0.7797291554114425
0.638907841781224   0.5431228030479904   0.7273950932858446   0.7478296085943323   0.5164192029922755   0.2419897750537278   0.7241924644954244   0.3173937398690268   0.5941382270565898   0.9115140115676151   0.8192047042882266   0.6275372669356836   0.9973787695960782   0.2689279559449034   0.4364503083297813   0.2891211329174514   0.07531308046905923   0.7173603511938136   0.8038643953503523   0.8239791252109   0.11853309677211   0.8709690424212279   0.2643246992612016   0.044249969799457466   0.47962525499088604   0.3278462393732374   0.536929605975357   0.2964203612051251   0.9632060519986105   0.08585646431950963   0.8127371414799326   0.9790266213360983   0.36906782494202073   0.17434245275189447   0.993532437191706   0.3514893544004148   0.37168905534594254   0.905414496806991   0.5570821288619248   0.06236822148296339   0.29637597487688333   0.18805414561317746   0.7532177335115725   0.2383890962720634   0.17784287810477334   0.3170851031919496   0.4888930342503709   0.19413912647260592   0.6982176231138872   0.9892388638187122   0.9519634282750139   0.8977187652674808   0.7350115711152767   0.9033823994992025   0.13922628679508128   0.9186921439313825   0.3659437461732559   0.7290399467473081   0.14569384960337525   0.5672027895309677   0.9942546908273133   0.823625449940317   0.5886117207414505   0.5048345680480043
0.69787871595043   0.6355713043271395   0.835393987229878   0.26644547177594097   0.5200358378456567   0.31848620113518994   0.3465009529795071   0.07230634530333503   0.8218182147317694   0.3292473373164777   0.39453752470449327   0.17458758003585423   0.08680664361649275   0.4258649378172752   0.25531123790941196   0.25589543610447174   0.7208628974432368   0.6968249910699671   0.10961738830603675   0.688692646573504   0.7266082066159235   0.8731995411296501   0.5210056675645862   0.18385807852549968   0.028729490665493462   0.23762823680251055   0.6856116803347082   0.9174126067495587   0.5086936528198368   0.9191420356673207   0.33911072735520104   0.8451062614462237   0.6868754380880674   0.5898946983508428   0.9445732026507078   0.6705186814103694   0.6000687944715746   0.16402976053356774   0.6892619647412958   0.4146232453058977   0.8792058970283377   0.4672047694636006   0.579644576435259   0.7259305987323937   0.15259769041241428   0.5940052283339505   0.05863890887067284   0.542072520206894   0.12386819974692083   0.35637699153144   0.37302722853596465   0.6246599134573353   0.6151745469270841   0.43723495586411937   0.0339165011807636   0.7795536520111116   0.9282991088390167   0.8473402575132765   0.0893432985300558   0.10903497060074213   0.3282303143674421   0.6833104969797087   0.40008133378876   0.6944117252948444
0.4490244173391043   0.2161057275161081   0.820436757353501   0.9684811265624507   0.29642672692669003   0.6221004991821575   0.761797848482828   0.42640860635555666   0.17255852717976922   0.26572350765071756   0.38877061994686346   0.8017486928982214   0.5573839802526852   0.8284885517865982   0.35485411876609985   0.0221950408871098   0.6290848714136685   0.9811482942733217   0.26551082023604405   0.9131600702863677   0.3008545570462264   0.297837797293613   0.865429486447284   0.21874834499152326   0.8518301397071221   0.08173206977750488   0.04499272909378309   0.25026721842907257   0.555403412780432   0.45963157059534737   0.283194880610955   0.8238586120735159   0.38284488560066277   0.1939080629446298   0.8944242606640915   0.022109919175294486   0.8254609053479776   0.3654195111580316   0.5395701418979917   0.9999148782881847   0.1963760339343091   0.38427121688470994   0.27405932166194763   0.08675480800181701   0.8955214768880827   0.08643341959109696   0.4086298352146636   0.8680064630102937   0.04369133718096068   0.004701349813592072   0.3636371061208805   0.6177392445812212   0.4882879244005287   0.5450697792182447   0.08044222550992552   0.7938806325077054   0.10544303879986593   0.3511617162736149   0.186017964845834   0.7717707133324108   0.2799821334518883   0.9857422051155833   0.6464478229478423   0.7718558350442262
0.08360609951757922   0.6014709882308733   0.3723885012858947   0.6851010270424092   0.1880846226294965   0.5150375686397763   0.9637586660712311   0.8170945640321153   0.1443932854485358   0.5103362188261843   0.6001215599503505   0.1993553194508942   0.6561053610480071   0.9652664396079396   0.519679334440425   0.4054746869431889   0.5506623222481412   0.6141047233343246   0.33366136959459103   0.633703973610778   0.2706801887962529   0.6283625182187415   0.6872135466467487   0.861848138566552   0.18707408927867364   0.026891529987868087   0.31482504536085404   0.17674711152414282   0.9989894666491772   0.5118539613480917   0.351066379289623   0.35965254749202746   0.8545961812006414   0.0015177425219074381   0.7509448193392725   0.16029722804113325   0.19849082015263422   0.036251302913967866   0.23126548489884743   0.7548225410979443   0.647828497904493   0.4221465795796432   0.8976041153042564   0.1211185674871663   0.37714830910824015   0.7937840613609018   0.2103905686575077   0.25927042892061436   0.19007421982956652   0.7668925313730337   0.8955655232966536   0.08252331739647156   0.19108475318038937   0.25503857002494196   0.5444991440070306   0.7228707699044441   0.336488571979748   0.25352082750303456   0.7935543246677582   0.5625735418633109   0.13799775182711377   0.21726952458906668   0.5622888397689108   0.8077510007653665
0.49016925392262073   0.7951229450094235   0.6646847244646543   0.6866324332782002   0.11302094481438059   0.001338883648521677   0.4542941558071467   0.4273620043575858   0.9229467249848141   0.23444635227548796   0.5587286325104931   0.34483868696111425   0.7318619718044247   0.979407782250546   0.014229488503462437   0.6219679170566701   0.39537339982467673   0.7258869547475114   0.22067516383570424   0.05939437519335928   0.25737564799756296   0.5086174301584447   0.6583863240667934   0.2516433744279928   0.7672063940749422   0.7134944851490213   0.9937015996021391   0.5650109411497926   0.6541854492605617   0.7121556015004996   0.5394074437949924   0.13764893679220677   0.7312387242757475   0.4777092492250117   0.9806788112844993   0.7928102498310925   0.9993767524713228   0.49830146697446565   0.9664493227810369   0.17084233277442235   0.6040033526466461   0.7724145122269542   0.7457741589453326   0.11144795758106307   0.34662770464908316   0.26379708206850944   0.08738783487853917   0.8598045831530703   0.5794213105741409   0.5503025969194881   0.09368623527640008   0.2947936420032777   0.9252358613135794   0.8381469954189885   0.5542787914814077   0.15714470521107093   0.1939971370378318   0.3604377461939769   0.5735999801969084   0.36433445537997844   0.194620384566509   0.8621362792195112   0.6071506574158715   0.1934921226055561
0.5906170319198629   0.089721766992557   0.8613764984705388   0.08204416502449302   0.24398932727077977   0.8259246849240476   0.7739886635919997   0.22223958187142273   0.6645680166966388   0.2756220880045594   0.6803024283155996   0.927445939868145   0.7393321553830594   0.4374750925855709   0.1260236368341919   0.7703012346570741   0.5453350183452277   0.07703734639159397   0.5524236566372835   0.4059667792770956   0.35071463377871864   0.21490106717208277   0.9452729992214121   0.21247465667153956   0.7600976018588557   0.12517930017952575   0.08389650075087328   0.13043049164704654   0.516108274588076   0.2992546152554782   0.30990783715887366   0.9081909097756238   0.8515402578914372   0.02363252725091882   0.6296054088432741   0.9807449699074787   0.11220810250837768   0.586157434665348   0.5035817720090822   0.2104437352504047   0.5668730841631501   0.509120088273754   0.9511581153717986   0.804476955973309   0.2161584503844314   0.29421902110167125   0.00588511615038655   0.5920022993017695   0.45606084852557566   0.16903972092214548   0.9219886153995133   0.461571807654723   0.9399525739374998   0.8697851056666672   0.6120807782406397   0.5533808978790992   0.08841231604606259   0.8461525784157484   0.9824753693973656   0.5726359279716204   0.9762042135376849   0.25999514375040045   0.4788935973882834   0.3621921927212157
0.40933112937453486   0.7508750554766465   0.5277354820164848   0.5577152367479067   0.19317267899010346   0.45665603437497526   0.5218503658660982   0.9657129374461372   0.7371118304645278   0.2876163134528298   0.599861750466585   0.5041411297914142   0.797159256527028   0.4178312077861625   0.9877809722259453   0.950760231912315   0.7087469404809654   0.5716786293704141   0.005305602828579719   0.3781243039406946   0.7325427269432806   0.31168348562001363   0.5264120054402963   0.01593211121947886   0.3232115975687457   0.5608084301433671   0.9986765234238116   0.45821687447157217   0.13003891857864222   0.10415239576839189   0.4768261575577134   0.492503937025435   0.3929270881141145   0.8165360823155621   0.8769644070911284   0.9883628072340208   0.5957678315870863   0.39870487452939957   0.8891834348651831   0.03760257532170579   0.8870208911061209   0.8270262451589855   0.8838778320366034   0.6594782713810112   0.15447816416284035   0.5153427595389719   0.3574658265963071   0.6435461601615323   0.8312665665940947   0.9545343293956048   0.3587893031724955   0.18532928568996015   0.7012276480154525   0.8503819336272128   0.8819631456147822   0.6928253486645252   0.308300559901338   0.03384585131165076   0.004998738523653685   0.7044625414305044   0.7125327283142516   0.6351409767822511   0.11581530365847051   0.6668599661087986
0.8255118372081307   0.8081147316232656   0.23193747162186704   0.007381694727787359   0.6710336730452903   0.2927719720842938   0.87447164502556   0.363835534566255   0.8397671064511957   0.33823764268868906   0.5156823418530644   0.17850624887629485   0.13853945843574325   0.4878557090614762   0.6337191962382822   0.4856809002117697   0.8302388985344052   0.4540098577498254   0.6287204577146286   0.7812183587812653   0.1177061702201537   0.8188688809675743   0.512905154056158   0.11435839267246677   0.292194333012023   0.010754149344308572   0.280967682434291   0.10697669794467941   0.6211606599667328   0.7179821772600148   0.4064960374087311   0.7431411633784244   0.7813935535155371   0.37974453457132573   0.8908136955556667   0.5646349145021295   0.6428540950797939   0.8918888255098496   0.2570944993173845   0.07895401429035985   0.8126151965453886   0.43787896776002416   0.6283740416027559   0.29773565550909453   0.6949090263252349   0.61901008679245   0.11546888754659791   0.18337726283662775   0.4027146933132118   0.6082559374481413   0.834501205112307   0.07640056489194834   0.7815540333464791   0.8902737601881265   0.42800516770357583   0.33325940151352396   0.00016047983094200904   0.5105292256168008   0.5371914721479092   0.7686244870113944   0.3573063847511482   0.6186404001069512   0.28009697283052465   0.6896704727210345
0.5446911882057596   0.18076143234692704   0.6517229312277687   0.39193481721194   0.8497821618805248   0.5617513455544771   0.5362540436811708   0.2085575543753123   0.44706746856731294   0.9534954081063357   0.7017528385688638   0.13215698948336393   0.6655134352208338   0.06322164791820914   0.273747670865288   0.79889758796984   0.6653529553898918   0.5526924223014084   0.7365561987173789   0.030273100958445577   0.30804657063874363   0.934052022194457   0.4564592258868542   0.340602628237411   0.7633553824329841   0.7532905898475301   0.8047362946590855   0.9486678110254709   0.9135732205524593   0.19153924429305294   0.2684822509779147   0.7401102566501587   0.4665057519851464   0.2380438361867172   0.5667294124090508   0.6079532671667948   0.8009923167643126   0.17482218826850807   0.29298174154376283   0.8090556791969548   0.1356393613744207   0.6221297659670998   0.5564255428263839   0.7787825782385092   0.827592790735677   0.6880777437726426   0.09996631693952972   0.43817995000109816   0.06423740830269302   0.9347871539251126   0.2952300222804442   0.4895121389756272   0.1506641877502337   0.7432479096320597   0.026747771302529463   0.7494018823254684   0.6841584357650874   0.5052040734453425   0.4600183588934786   0.14144861515867374   0.8831661190007748   0.3303818851768344   0.16703661734971575   0.332392935961719
0.7475267576263541   0.7082521192097346   0.6106110745233319   0.5536103577232098   0.9199339668906771   0.020174375437092013   0.5106447575838021   0.1154304077221116   0.855696558587984   0.0853872215119794   0.2154147353033579   0.6259182687464844   0.7050323708377503   0.34213931187991975   0.1886669640008284   0.8765163864210159   0.020873935072662955   0.8369352384345773   0.7286486051073499   0.7350677712623422   0.13770781607188814   0.5065533532577429   0.5616119877576341   0.4026748353006232   0.3901810584455341   0.7983012340480082   0.9510009132343022   0.8490644775774134   0.47024709155485706   0.7781268586109161   0.4403561556505002   0.7336340698553019   0.614550532966873   0.6927396370989368   0.2249414203471423   0.10771580110881744   0.9095181621291227   0.3506003252190171   0.036274456346313856   0.23119941468780153   0.8886442270564597   0.5136650867844398   0.307625851238964   0.49613164342545935   0.7509364109845716   0.007111733526696943   0.7460138634813299   0.09345680812483612   0.36075535253903757   0.20881049947868877   0.7950129502470277   0.24439233054742265   0.8905082609841806   0.4306836408677726   0.35465679459652755   0.5107582606921208   0.2759577280173075   0.7379440037688358   0.12971537424938526   0.40304245958330337   0.3664395658881847   0.38734367854981877   0.09344091790307141   0.17184304489550184
0.4777953388317249   0.873678591765379   0.7858150666641074   0.6757114014700425   0.7268589278471533   0.8665668582386821   0.039801203182777405   0.5822545933452064   0.36610357530811577   0.6577563587599933   0.24478825293574968   0.33786226279778375   0.47559531432393526   0.2270727178922207   0.8901314583392221   0.8271040021056629   0.19963758630662776   0.4891287141233849   0.7604160840898369   0.42406154252235956   0.833198020418443   0.10178503557356611   0.6669751661867654   0.2522184976268578   0.35540268158671806   0.22810644380818715   0.8811600995226581   0.5765070961568153   0.6285437537395647   0.3615395855695051   0.8413588963398807   0.9942525028116088   0.262440178431449   0.7037832268095119   0.596570643404131   0.6563902400138252   0.7868448641075138   0.47671050891729116   0.7064391850649089   0.8292862379081622   0.587207277800886   0.9875817947939063   0.946023100975072   0.40522469538580264   0.754009257382443   0.8857967592203402   0.2790479347883065   0.1530061977589449   0.3986065757957249   0.6576903154121531   0.3978878352656484   0.5764991016021296   0.7700628220561602   0.29615072984264795   0.5565289389257677   0.5822465987905208   0.5076226436247111   0.5923675030331361   0.9599582955216367   0.9258563587766956   0.7207777795171973   0.11565699411584493   0.2535191104567278   0.09657012086853342
0.13357050171631135   0.12807519932193864   0.30749600948165584   0.6913454254827308   0.37956124433386834   0.24227844010159846   0.028448074693349354   0.538339227723786   0.9809546685381435   0.5845881246894454   0.630560239427701   0.9618401261216563   0.2108918464819833   0.2884373948467975   0.07403130050193327   0.37959352733113555   0.7032692028572722   0.6960698918136614   0.11407300498029659   0.4537371685544399   0.9824914233400748   0.5804128976978165   0.8605538945235688   0.35716704768590646   0.8489209216237634   0.45233769837587784   0.5530578850419129   0.6658216222031756   0.4693596772898951   0.21005925827427938   0.5246098103485636   0.12748239447938978   0.48840500875175163   0.625471133584834   0.8940495709208626   0.1656422683577335   0.2775131622697683   0.3370337387380365   0.8200182704189294   0.7860487410265979   0.5742439594124962   0.640963846924375   0.7059452654386328   0.3323115724721581   0.5917525360724213   0.06055094922655862   0.845391370915064   0.9751445247862516   0.7428316144486579   0.6082132508506808   0.29233348587315106   0.3093229025830759   0.2734719371587627   0.39815399257640144   0.7677236755245875   0.1818405081036861   0.7850669284070111   0.7726828589915675   0.8736741046037249   0.01619823974595261   0.5075537661372428   0.43564912025353103   0.05365583418479554   0.23014949871935464
0.9333098067247466   0.794685273329156   0.3477105687461628   0.8978379262471966   0.34155727065232533   0.7341343241025973   0.5023191978310988   0.9226934014609449   0.5987256562036675   0.1259210732519165   0.20998571195794777   0.6133704988778691   0.32525371904490474   0.7277670806755151   0.44226203643336026   0.43152999077418297   0.5401867906378937   0.9550842216839476   0.5685879318296354   0.41533175102823033   0.03263302450065085   0.5194351014304166   0.5149320976448398   0.18518225230887572   0.09932321777590422   0.7247498281012607   0.16722152889867709   0.28734432606167915   0.7577659471235789   0.9906155039986634   0.6649023310675782   0.3646509246007342   0.15904029091991143   0.8646944307467468   0.4549166191096305   0.7512804257228651   0.8337865718750067   0.13692735007123172   0.012654582676270202   0.31975043494868216   0.29359978123711306   0.18184312838728411   0.44406665084663477   0.9044186839204518   0.2609667567364622   0.6624080269568675   0.9291345532017949   0.7192364316115761   0.161643538960558   0.9376581988556069   0.7619130243031178   0.43189210554989693   0.40387759183697913   0.9470426948569436   0.09701069323553957   0.06724118094916272   0.24483730091706768   0.08234826411019676   0.6420940741259091   0.3159607552262976   0.41105072904206097   0.945420914038965   0.6294394914496388   0.9962103202776154
0.11745094780494791   0.7635777856516809   0.1853728406030041   0.09179163635716359   0.8564841910684857   0.10116975869481337   0.2562382874012092   0.3725552047455875   0.6948406521079277   0.16351155983920648   0.4943252630980913   0.9406630991956906   0.2909630602709486   0.2164688649822629   0.39731456986255176   0.8734219182465278   0.046125759353880906   0.13412060087206615   0.7552204957366427   0.5574611630202303   0.6350750303118199   0.18869968683310112   0.1257810042870038   0.5612508427426148   0.517624082506872   0.4251219011814202   0.9404081636839997   0.46945920638545124   0.6611398914383864   0.32395214248660686   0.6841698762827906   0.09690400163986378   0.9662992393304586   0.16044058264740038   0.18984461318469917   0.1562409024441732   0.67533617905951   0.9439717176651374   0.7925300433221474   0.28281898419764534   0.6292104197056291   0.8098511167930713   0.03730954758550471   0.7253578211774151   0.9941353893938092   0.6211514299599702   0.9115285432985009   0.1641069784348002   0.4765113068869372   0.19602952877854998   0.9711203796145012   0.6946477720493489   0.8153714154485509   0.8720773862919432   0.2869505033317107   0.5977437704094852   0.8490721761180923   0.7116368036445427   0.09710589014701149   0.44150286796531196   0.17373599705858225   0.7676650859794053   0.30457584682486405   0.15868388376766662
0.5445255773529531   0.957813969186334   0.26726629923935935   0.4333260625902515   0.550390187959144   0.3366625392263638   0.35573775594085844   0.2692190841554513   0.07387888107220673   0.1406330104478138   0.3846173763263573   0.5745713121061023   0.25850746562365584   0.26855562415587064   0.0976668729946466   0.9768275416966172   0.40943528950556357   0.5569188205113279   0.0005609828476351168   0.5353246737313052   0.23569929244698135   0.7892537345319226   0.695985136022771   0.3766407899636386   0.6911737150940283   0.8314397653455886   0.42871883678341166   0.9433147273733871   0.1407835271348843   0.49477722611922476   0.07298108084255323   0.6740956432179357   0.06690464606267756   0.35414421567141097   0.688363704516196   0.09952433111183331   0.8083971804390218   0.08558859151554034   0.5906968315215494   0.12269678941521613   0.39896189093345813   0.5286697710042124   0.5901358486739142   0.5873721156839109   0.16326259848647678   0.7394160364722899   0.8941507126511432   0.21073132572027237   0.47208888339244853   0.9079762711267013   0.46543187586773155   0.26741659834688536   0.33130535625756424   0.4131990450074766   0.3924507950251783   0.5933209551289497   0.2644007101948867   0.05905482933606562   0.7040870905089823   0.4937966240171163   0.456003529755865   0.9734662378205253   0.11339025898743296   0.3710998346019002
0.05704163882240687   0.4447964668163128   0.5232544103135187   0.7837277189179893   0.8937790403359301   0.7053804303440229   0.6291036976623755   0.5729963931977169   0.42169015694348155   0.7974041592173216   0.16367182179464398   0.3055797948508316   0.09038480068591728   0.38420511420984493   0.7712210267694657   0.712258839721882   0.8259840904910306   0.3251502848737793   0.06713393626048335   0.2184622157047656   0.3699805607351656   0.351684047053254   0.9537436772730504   0.8473623811028654   0.31293892191275874   0.9068875802369412   0.43048926695953166   0.06363466218487611   0.41915988157682865   0.2015071498929183   0.8013855692971561   0.4906382689871592   0.997469724633347   0.4041029906755968   0.6377137475025122   0.18505847413632756   0.9070849239474298   0.01989787646575184   0.8664927207330465   0.4727996344144456   0.08110083345639922   0.6947475915919725   0.7993587844725631   0.25433741870968   0.7111202727212337   0.3430635445387185   0.8456151071995127   0.40697503760681464   0.39818135080847494   0.43617596430177735   0.4151258402399811   0.3433403754219385   0.9790214692316463   0.23466881440885903   0.613740270942825   0.8527021064347794   0.9815517445982992   0.8305658237332623   0.9760265234403128   0.6676436322984518   0.0744668206508694   0.8106679472675105   0.10953380270726631   0.19484399788400614
0.9933659871944702   0.11592035567553789   0.31017501823470317   0.9405065791743261   0.28224571447323654   0.7728568111368194   0.4645599110351904   0.5335315415675115   0.8840643636647616   0.336680846835042   0.049434070795209305   0.19019116614557297   0.9050428944331154   0.10201203242618298   0.4356937998523843   0.3374890597107936   0.9234911498348161   0.2714462086929207   0.45966727641207156   0.6698454274123419   0.8490243291839467   0.4607782614254103   0.35013347370480524   0.4750014295283357   0.8556583419894765   0.3448579057498724   0.039958455470102044   0.5344948503540096   0.57341262751624   0.572001094613053   0.5753985444349117   0.0009633087864980596   0.6893482638514784   0.235320247778011   0.5259644736397023   0.8107721426409251   0.784305369418363   0.13330821535182802   0.09027067378731798   0.4732830829301315   0.860814219583547   0.8618620066589073   0.6306033973752464   0.8034376555177897   0.01178989039960025   0.40108374523349705   0.2804699236704412   0.328436225989454   0.15613154841012372   0.056225839483624675   0.2405114682003392   0.7939413756354444   0.5827189208938837   0.48422474487057166   0.6651129237654275   0.7929780668489463   0.8933706570424054   0.24890449709256066   0.13914845012572524   0.9822059242080212   0.10906528762404225   0.11559628174073261   0.048877776338407244   0.5089228412778898
0.2482510680404953   0.2537342750818253   0.4182743789631608   0.7054851857601001   0.23646117764089505   0.8526505298483282   0.13780445529271956   0.3770489597706462   0.08032962923077133   0.7964246903647035   0.8972929870923804   0.5831075841352017   0.49761070833688764   0.3121999454941319   0.23218006332695282   0.7901295172862554   0.6042400512944823   0.06329544840157127   0.0930316132012276   0.8079235930782341   0.49517476367044005   0.9476991666608386   0.04415383686282035   0.2990007518003443   0.24692369562994476   0.6939648915790133   0.6258794578996596   0.5935155660402441   0.010462517989049711   0.8413143617306851   0.48807500260694   0.21646660626959802   0.9301328887582784   0.04488967136598157   0.5907820155145596   0.6333590221343963   0.43252218042139073   0.7326897258718497   0.35860195218760677   0.843229504848141   0.8282821291269085   0.6693942774702784   0.26557033898637916   0.035305911769906835   0.3331073654564684   0.7216951108094397   0.22141650212355884   0.7363051599695626   0.08618366982652366   0.027730219230426394   0.5955370442238993   0.14278959392931836   0.07572115183747394   0.18641585749974127   0.10746204161695928   0.9263229876597203   0.14558826307919556   0.1415261861337597   0.5166800261023997   0.29296396552532405   0.7130660826578048   0.40883646026191   0.1580780739147929   0.44973446067718315
0.8847839535308963   0.7394421827916317   0.8925077349284137   0.4144285489072763   0.551676588074428   0.01774707198219187   0.6710912328048548   0.6781233889377137   0.4654929182479043   0.9900168527517654   0.07555418858095561   0.5353337950083954   0.3897717664104303   0.8036009952520242   0.9680921469639964   0.6090108073486751   0.24418350333123479   0.6620748091182646   0.45141212086159666   0.316046841823351   0.5311174206734299   0.2532383488563545   0.29333404694680376   0.8663123811461678   0.6463334671425336   0.5137961660647229   0.40082631201839003   0.45188383223889156   0.0946568790681057   0.496049094082531   0.7297350792135352   0.7737604433011778   0.6291639608202014   0.5060322413307655   0.6541808906325796   0.23842664829278237   0.23939219440977108   0.7024312460787413   0.6860887436685832   0.6294158409441073   0.9952086910785363   0.0403564369604768   0.23467662280698656   0.31336899912075633   0.46409127040510634   0.7871180881041223   0.9413425758601828   0.44705661797458845   0.8177578032625726   0.2733219220393994   0.5405162638417927   0.9951727857356969   0.723100924194467   0.7772728279568685   0.8107811846282577   0.2214123424345191   0.09393696337426556   0.2712405866261029   0.1566002939956781   0.9829856941417368   0.8545447689644945   0.5688093405473617   0.4705115503270949   0.3535698531976294
0.8593360778859582   0.5284529035868848   0.23583492752010835   0.04020085407687307   0.3952448074808519   0.7413348154827625   0.2944923516599255   0.5931442361022846   0.5774870042182791   0.46801289344336305   0.7539760878181327   0.5979714503665877   0.8543860800238122   0.6907400654864946   0.9431949031898751   0.37655910793206865   0.7604491166495466   0.4194994788603917   0.786594609194197   0.39357341379033195   0.9059043476850521   0.8506901383130301   0.3160830588671021   0.04000356059270255   0.046568269799093974   0.3222372347261453   0.08024813134699375   0.9998027065158295   0.6513234623182421   0.5809024192433828   0.7857557796870682   0.40665847041354486   0.07383645809996292   0.11288952580001974   0.031779691868935506   0.8086870200469571   0.21945037807615073   0.4221494603135251   0.08858478867906043   0.4321279121148885   0.4590012614266041   0.002649981453133424   0.30199017948486345   0.038554498324556534   0.5530969137415519   0.15195984314010333   0.9859071206177613   0.998550937731854   0.5065286439424579   0.8297226084139581   0.9056589892707676   0.9987482312160245   0.8552051816242159   0.24882018917057527   0.11990320958369938   0.5920897608024797   0.7813687235242529   0.13593066337055554   0.08812351771476387   0.7834027407555225   0.5619183454481022   0.7137812030570304   0.9995387290357034   0.3512748286406341
0.10291708402149813   0.711131221603897   0.69754854955084   0.31272033031607754   0.5498201702799462   0.5591713784637936   0.7116414289330787   0.31416939258422355   0.043291526337488284   0.7294487700498355   0.805982439662311   0.31542116136819903   0.18808634471327246   0.48062858087926036   0.6860792300786116   0.7233314005657194   0.40671762118901955   0.3446979175087048   0.5979557123638478   0.9399286598101968   0.8447992757409173   0.6309167144516744   0.5984169833281443   0.5886538311695627   0.7418821917194192   0.9197854928477774   0.9008684337773043   0.27593350085348517   0.19206202143947299   0.3606141143839838   0.18922700484422567   0.9617641082692616   0.1487704951019847   0.6311653443341482   0.38324456518191463   0.6463429469010625   0.9606841503887122   0.1505367634548878   0.697165335103303   0.9230115463353432   0.5539665291996927   0.805838845946183   0.09920962273945524   0.9830828865251463   0.7091672534587754   0.1749221314945086   0.5007926394113109   0.3944290553555836   0.9672850617393561   0.2551366386467312   0.5999242056340066   0.11849555450209838   0.7752230402998832   0.8945225242627474   0.41069720078978095   0.15673144623283675   0.6264525451978985   0.26335717992859925   0.02745263560786631   0.5103884993317742   0.6657683948091863   0.11282041647371142   0.3302873005045633   0.587376952996431
0.1118018656094935   0.30698157052752845   0.23107767776510804   0.6042940664712847   0.4026346121507181   0.1320594390330198   0.7302850383537971   0.2098650111157011   0.4353495504113619   0.8769228003862887   0.1303608327197905   0.09136945661360271   0.6601265101114787   0.9824002761235412   0.7196636319300095   0.934638010380766   0.03367396491358027   0.719043096194942   0.6922109963221432   0.4242495110489918   0.36790557010439406   0.6062226797212306   0.36192369581757994   0.8368725580525608   0.25610370449490055   0.2992411091937021   0.13084601805247187   0.23257849158127608   0.8534690923441824   0.1671816701606823   0.40056097969867477   0.022713480465574972   0.4181195419328205   0.2902588697743937   0.2702001469788843   0.9313440238519722   0.7579930318213418   0.30785859365085244   0.5505365150488748   0.9967060134712062   0.7243190669077615   0.5888154974559104   0.8583255187267316   0.5724565024222146   0.3564134968033674   0.9825928177346799   0.49640182290915164   0.7355839443696538   0.10030979230846689   0.6833517085409778   0.36555580485667977   0.5030054527883777   0.24684069996428445   0.5161700383802955   0.964994825158005   0.48029197232280274   0.828721158031464   0.22591116860590182   0.6947946781791208   0.5489479484708305   0.07072812621012217   0.9180525749550493   0.14425816313024595   0.5522419349996242
0.34640905930236066   0.3292370774991389   0.2859326444035144   0.9797854325774097   0.9899955624989932   0.346644259764459   0.7895308214943627   0.24420148820775586   0.8896857701905263   0.6632925512234812   0.42397501663768294   0.7411960354193782   0.6428450702262419   0.14712251284318573   0.45898019147967795   0.26090406309657543   0.814123912194778   0.9212113442372839   0.7641855133005572   0.7119561146257449   0.7433957859846558   0.0031587692822345323   0.6199273501703112   0.15971417962612078   0.3969867266822951   0.6739216917830956   0.33399470576679685   0.17992874704871115   0.4069911641833019   0.3272774320186366   0.5444638842724341   0.9357272588409553   0.5173053939927755   0.6639848807951554   0.12048886763475114   0.19453122342157708   0.8744603237665336   0.5168623679519697   0.6615086761550732   0.9336271603250017   0.060336411571755635   0.5956510237146858   0.897323162854516   0.2216710456992567   0.31694062558709984   0.5924922544324512   0.2773958126842047   0.06195686607313591   0.9199538989048047   0.9185705626493557   0.9434011069174079   0.8820281190244248   0.5129627347215028   0.591293130630719   0.3989372226449738   0.9463008601834695   0.9956573407287272   0.9273082498355636   0.27844835501022264   0.7517696367618925   0.12119701696219366   0.4104458818835939   0.6169396788551494   0.8181424764368908
0.06086060539043803   0.8147948581689081   0.7196165160006335   0.5964714307376341   0.7439199798033382   0.22230260373645686   0.4422207033164287   0.5345145646644982   0.8239660808985335   0.3037320410871012   0.49881959639902085   0.6524864456400734   0.3110033461770307   0.7124389104563822   0.09988237375404707   0.7061855854566038   0.31534600544830343   0.7851306606208186   0.8214340187438245   0.9544159486947115   0.19414898848610979   0.3746847787372247   0.20449433988867502   0.13627347225782066   0.13328838309567176   0.5598899205683167   0.48487782388804157   0.5398020415201866   0.3893684032923335   0.3375873168318598   0.04265712057161285   0.005287476855688447   0.5654023223938001   0.033855275744758564   0.543837524172592   0.35280103121561507   0.2543989762167693   0.32141636528837636   0.44395515041854494   0.6466154457590112   0.9390529707684658   0.5362857046675578   0.6225211316747205   0.6921994970642997   0.7449039822823561   0.161600925930333   0.41802679178604546   0.5559260248064791   0.6116155991866844   0.6017110053620164   0.933148967898004   0.016123983286292512   0.22224719589435082   0.2641236885301566   0.8904918473263911   0.010836506430604066   0.6568448735005508   0.23026841278539806   0.34665432315379907   0.658035475214989   0.4024458972837815   0.9088520474970216   0.9026991727352541   0.011420029455977775
0.4633929265153156   0.37256634282946394   0.2801780410605336   0.31922053239167797   0.7184889442329595   0.21096541689913093   0.8621512492744882   0.7632945075851989   0.10687334504627512   0.6092544115371146   0.9290022813764842   0.7471705242989064   0.8846261491519243   0.3451307230069579   0.03851043405009317   0.7363340178683023   0.22778127565137352   0.11486231022155984   0.6918561108962941   0.0782985426533133   0.8253353783675921   0.20601026272453815   0.78915693816104   0.06687851319733554   0.36194245185227647   0.8334439198950742   0.5089788971005064   0.7476579808056575   0.643453507619317   0.6224785029959433   0.6468276478260182   0.9843634732204587   0.5365801625730419   0.013224091458828762   0.717825366449534   0.2371929489215523   0.6519540134211176   0.6680933684518708   0.6793149323994409   0.50085893105325   0.42417273776974407   0.553231058230311   0.9874588215031467   0.4225603883999367   0.598837359402152   0.3472207955057729   0.19830188334210672   0.35568187520260114   0.23689490754987558   0.5137768756106986   0.6893229862416004   0.6080238943969436   0.5934413999305586   0.8912983726147554   0.0424953384155821   0.6236604211764849   0.056861237357516733   0.8780742811559267   0.3246699719660481   0.38646747225493266   0.40490722393639916   0.20998091270405575   0.6453550395666072   0.8856085412016826
0.980734486166655   0.6567498544737448   0.6578962180634605   0.463048152801746   0.38189712676450305   0.3095290589679719   0.4595943347213538   0.10736627759914483   0.14500221921462747   0.7957521833572732   0.7702713484797534   0.4993423832022012   0.5515608192840689   0.9044538107425178   0.7277760100641714   0.8756819620257162   0.4946995819265521   0.026379529586591188   0.4031060380981233   0.4892144897707836   0.08979235799015298   0.8163986168825355   0.7577509985315161   0.6036059485691009   0.1090578718234979   0.1596487624087907   0.09985478046805552   0.14055779576735494   0.7271607450589949   0.8501197034408188   0.6402604457467017   0.03319151816821012   0.5821585258443673   0.05436752008354562   0.8699890972669483   0.5338491349660089   0.0305977065602985   0.1499137093410278   0.14221308720277692   0.6581671729402927   0.5358981246337463   0.12353417975443662   0.7391070491046536   0.16895268316950907   0.44610576664359336   0.3071355628719012   0.9813560505731377   0.5653467346004082   0.3370478948200955   0.1474868004631105   0.8815012701050822   0.4247889388330532   0.6098871497611006   0.2973670970222917   0.24124082435838037   0.39159742066484304   0.02772862391673327   0.24299957693874608   0.3712517270914321   0.8577482856988341   0.9971309173564348   0.09308586759771827   0.22903863988865517   0.19958111275854148
0.4612327927226884   0.9695516878432816   0.4899315907840015   0.030628429589032422   0.015127026079095027   0.6624161249713805   0.5085755402108639   0.46528169498862426   0.6780791312589995   0.51492932450827   0.6270742701057818   0.04049275615557108   0.0681919814978989   0.21756222748597825   0.38583344574740136   0.648895335490728   0.04046335758116563   0.9745626505472322   0.014581718655969269   0.7911470497918939   0.04333244022473086   0.8814767829495139   0.7855430787673141   0.5915659370333524   0.5820996475020425   0.9119250951062323   0.2956114879833126   0.5609375074443199   0.5669726214229475   0.24950897013485182   0.7870359477724487   0.09565581245569567   0.8888934901639479   0.7345796456265818   0.15996167766666694   0.05516305630012459   0.820701508666049   0.5170174181406036   0.7741282319192656   0.40626772080939655   0.7802381510848834   0.5424547675933714   0.7595465132632963   0.6151206710175027   0.7369057108601524   0.6609779846438575   0.9740034344959823   0.023554733984150346   0.15480606335811004   0.7490528895376252   0.6783919465126697   0.4626172265398304   0.5878334419351626   0.4995439194027734   0.8913559987402209   0.36696141408413474   0.6989399517712147   0.7649642737761915   0.731394321073554   0.31179835778401016   0.8782384431051657   0.24794685563558788   0.9572660891542885   0.9055306369746136
0.09800029202028242   0.7054920880422165   0.19771957589099212   0.2904099659571108   0.36109458116012993   0.04451410339835899   0.22371614139500992   0.2668552319729605   0.20628851780201987   0.29546121386073376   0.5453241948823403   0.8042380054331301   0.6184550758668572   0.7959172944579604   0.6539681961421194   0.4372765913489954   0.9195151240956425   0.030953020681768913   0.9225738750685654   0.12547823356498525   0.04127668099047674   0.783006165046181   0.965307785914277   0.21994759659037166   0.9432763889701943   0.07751407700396455   0.7675882100232849   0.9295376306332608   0.5821818078100645   0.03299997360560556   0.543872068628275   0.6626823986603003   0.37589329000804456   0.7375387597448718   0.9985478737459347   0.8584443932271701   0.7574382141411873   0.9416214652869114   0.3445796776038153   0.4211678018781748   0.8379230900455448   0.9106684446051424   0.4220058025352499   0.2956895683131896   0.796646409055068   0.12766227955896142   0.4566980166209729   0.07574197172281791   0.8533700200848737   0.05014820255499687   0.6891098065976881   0.14620434108955707   0.27118821227480927   0.01714822894939131   0.14523773796941306   0.4835219424292568   0.8952949222667648   0.2796094692045195   0.1466898642234784   0.6250775492020866   0.1378567081255775   0.3379880039176082   0.8021101866196632   0.20390974732391176
0.2999336180800327   0.42731955931246574   0.3801043840844132   0.9082201790107222   0.5032872090249647   0.2996572797535043   0.9234063674634403   0.8324782072879043   0.649917188940091   0.24950907719850746   0.2342965608657523   0.6862738661983472   0.37872897666528166   0.23236084824911613   0.08905882289633922   0.20275192376909043   0.4834340543985169   0.9527513790445966   0.9423689586728609   0.5776743745670039   0.3455773462729394   0.6147633751269884   0.1402587720531977   0.37376462724309206   0.04564372819290671   0.18744381581452269   0.7601543879687845   0.4655444482323699   0.542356519167942   0.8877865360610183   0.8367480205053441   0.6330662409444656   0.892439330227851   0.6382774588625109   0.6024514596395919   0.9467923747461184   0.5137103535625693   0.4059166106133948   0.5133926367432526   0.744040450977028   0.03027629916405245   0.4531652315687982   0.5710236780703918   0.16636607641002413   0.684698952891113   0.8384018564418098   0.4307649060171941   0.7926014491669321   0.6390552246982063   0.6509580406272871   0.6706105180484097   0.32705700093456214   0.09669870553026429   0.7631715045662687   0.8338624975430654   0.6939907599900965   0.20425937530241325   0.12489404570375781   0.2314110379034736   0.7471983852439782   0.6905490217398439   0.718977435090363   0.718018401160221   0.0031579342669501606
0.6602727225757914   0.26581220352156487   0.14699472308982914   0.836791857856926   0.9755737696846785   0.42741034707975506   0.716229817072635   0.04419040868999397   0.3365185449864721   0.776452306452468   0.0456192990242254   0.7171334077554318   0.2398198394562078   0.013280801886199265   0.21175680148115994   0.02314264776533526   0.03556046415379456   0.8883867561824415   0.9803457635776863   0.2759442625213571   0.34501144241395065   0.1694093210920784   0.2623273624174654   0.27278632825440696   0.6847387198381593   0.9035971175705135   0.11533263932763628   0.4359944703974809   0.7091649501534808   0.47618677049075847   0.39910282225500127   0.39180406170748694   0.37264640516700875   0.6997344640382904   0.35348352323077586   0.6746706539520552   0.13282656571080095   0.6864536621520912   0.1417267217496159   0.6515280061867199   0.09726610155700639   0.7980669059696498   0.16138095817192954   0.3755837436653628   0.7522546591430557   0.6286575848775714   0.8990535957544641   0.10279741541095583   0.06751593930489647   0.7250604673070578   0.7837209564268278   0.6668029450134749   0.3583509891514156   0.2488736968162993   0.3846181341718266   0.27499888330598793   0.9857045839844069   0.5491392327780088   0.031134610941050758   0.6003282293539328   0.8528780182736059   0.8626855706259177   0.8894078891914349   0.9488002231672129
0.7556119167165996   0.06461866465626788   0.7280269310195053   0.5732164795018501   0.0033572575735438042   0.4359610797786965   0.8289733352650411   0.4704190640908943   0.9358413182686474   0.7109006124716387   0.04525237883821332   0.8036161190774194   0.5774903291172317   0.46202691565533943   0.6606342446663868   0.5286172357714315   0.5917857451328249   0.9128876828773306   0.6294996337253359   0.9282890064174987   0.738907726859219   0.05020211225141293   0.7400917445339011   0.9794887832502858   0.9832958101426195   0.985583447595145   0.012064813514395787   0.40627230374843565   0.9799385525690757   0.5496223678164486   0.18309147824935462   0.9358532396575414   0.0440972343004283   0.8387217553448097   0.13783909941114128   0.132237120580122   0.4666069051831966   0.3766948396894704   0.4772048547447546   0.6036198848086906   0.8748211600503717   0.4638071568121398   0.8477052210194186   0.6753308783911919   0.13591343319115273   0.4136050445607269   0.10761347648551753   0.6958420951409061   0.15261762304853327   0.42802159696558184   0.09554866297112173   0.2895697913924704   0.17267907047945763   0.8783992291491333   0.9124571847217672   0.353716551734929   0.12858183617902932   0.03967747380432351   0.7746180853106258   0.22147943115480703   0.6619749309958327   0.6629826341148531   0.29741323056587127   0.6178595463461165
0.787153770945461   0.19917547730271332   0.4497080095464526   0.9425286679549246   0.6512403377543083   0.7855704327419865   0.3420945330609351   0.24668657281401857   0.49862271470577507   0.35754883577640456   0.24654587008981338   0.9571167814215482   0.32594364422631744   0.4791496066272713   0.33408868536804626   0.6034002296866191   0.1973618080472881   0.4394721328229478   0.5594706000574204   0.3819207985318121   0.5353868770514554   0.7764894987080947   0.2620573694915492   0.7640612521856956   0.7482331061059943   0.5773140214053814   0.8123493599450965   0.821532584230771   0.09699276835168592   0.7917435886633949   0.4702548268841614   0.5748460114167524   0.5983700536459109   0.43419475288699033   0.22370895679434807   0.6177292299952043   0.27242640941959345   0.955045146259719   0.8896202714263018   0.014329000308585142   0.07506460137230535   0.5155730134367713   0.3301496713688814   0.632408201776773   0.53967772432085   0.7390835147286766   0.06809230187733224   0.8683469495910774   0.7914446182148558   0.16176949332329532   0.25574294193223573   0.046814365360306365   0.6944518498631698   0.37002590465990043   0.7854881150480743   0.4719683539435539   0.09608179621725894   0.9358311517729101   0.5617791582537263   0.8542391239483497   0.8236553867976655   0.9807860055131911   0.6721588868274244   0.8399101236397645
0.7485907854253602   0.46521299207641975   0.342009215458543   0.20750192186299146   0.20891306110451013   0.7261294773477431   0.27391691358121073   0.3391549722719141   0.4174684428896544   0.5643599840244478   0.01817397164897504   0.29234060691160774   0.7230165930264846   0.19433407936454739   0.23268585660090074   0.8203722529680538   0.6269347968092256   0.2585029275916373   0.6709066983471745   0.9661331290197042   0.8032794100115601   0.2777169220784463   0.9987478115197501   0.12622300537993972   0.05468862458619996   0.8125039300020266   0.6567385960612071   0.9187210835169483   0.8457755634816898   0.08637445265428344   0.3828216824799964   0.5795661112450341   0.42830712059203546   0.5220144686298357   0.3646477108310213   0.2872255043334264   0.7052905275655509   0.3276803892652883   0.13196185423012058   0.4668532513653726   0.07835573075632525   0.06917746167365099   0.46105515588294604   0.5007201223456684   0.2750763207447651   0.7914605395952047   0.4623073443631959   0.3744971169657287   0.22038769615856518   0.9789566095931782   0.8055687483019888   0.4557760334487805   0.3746121326768753   0.8925821569388948   0.42274706582199245   0.8762099222037463   0.9463050120848399   0.37056768830905906   0.0580993549909711   0.5889844178703199   0.24101448451928903   0.04288729904377078   0.9261375007608506   0.12213116650494729
0.1626587537629638   0.9737098373701198   0.4650823448779045   0.6214110441592788   0.8875824330181986   0.18224929777491508   0.002775000514708561   0.24691392719355018   0.6671947368596335   0.20329268818173693   0.19720625221271976   0.7911378937447697   0.2925826041827581   0.3107105312428422   0.7744591863907273   0.9149279715410235   0.34627759209791825   0.9401428429337831   0.7163598313997562   0.32594355367070355   0.1052631075786292   0.8972555438900123   0.7902223306389057   0.20381238716575623   0.9426043538156654   0.9235457065198925   0.3251399857610012   0.5824013430064774   0.05502192079746677   0.7412964087449775   0.32236498524629265   0.3354874158129272   0.3878271839378333   0.5380037205632405   0.1251587330335729   0.5443495220681575   0.09524457975507515   0.22729318932039833   0.3506995466428456   0.629421550527134   0.748966987657157   0.28715034638661524   0.6343397152430893   0.3034779968564305   0.6437038800785277   0.3898948024966029   0.8441173846041836   0.09966560969067428   0.7010995262628623   0.46634909597671037   0.5189773988431824   0.5172642666841969   0.6460776054653955   0.7250526872317329   0.19661241359688975   0.18177685087126977   0.2582504215275622   0.1870489666684924   0.07145368056331684   0.6374273288031124   0.1630058417724871   0.959755777348094   0.7207541339204713   0.008005778275978297
0.4140388541153302   0.6726054309614788   0.08641441867738194   0.7045277814195477   0.7703349740368025   0.282710628464876   0.2422970340731983   0.6048621717288735   0.06923544777394015   0.8163615324881656   0.7233196352300159   0.08759790504467654   0.42315784230854464   0.09130884525643267   0.5267072216331261   0.9058210541734067   0.1649074207809824   0.9042598785879402   0.4552535410698093   0.26839372537029443   0.001901579008495279   0.9445041012398462   0.734499407149338   0.2603879470943161   0.587862724893165   0.27189867027836734   0.6480849884719562   0.5558601656747684   0.8175277508563626   0.9891880418134914   0.4057879543987578   0.9509979939458949   0.7482923030824224   0.17282650932532576   0.682468319168742   0.8634000889012183   0.32513446077387786   0.08151766406889308   0.15576109753561573   0.9575790347278116   0.16022703999289548   0.1772577854809528   0.7005075564658064   0.6891853093575171   0.1583254609844002   0.23275368424110662   0.9660081493164684   0.428797362263201   0.5704627360912351   0.9608550139627393   0.3179231608445122   0.8729371965884326   0.7529349852348725   0.971666972149248   0.9121352064457544   0.9219392026425377   0.004642682152449981   0.7988404628239222   0.22966688727701254   0.058539113741319405   0.6795082213785721   0.7173227987550291   0.07390578974139679   0.10096007901350786
0.5192811813856766   0.5400650132740763   0.37339823327559035   0.41177476965599075   0.36095572040127644   0.3073113290329697   0.407390083959122   0.9829774073927898   0.7904929843100413   0.3464563150702304   0.08946692311460977   0.1100402108043572   0.037557999075168866   0.3747893429209824   0.17733171666885533   0.1881010081618195   0.03291531692271888   0.5759488800970602   0.9476648293918428   0.1295618944205001   0.3534070955441468   0.858626081342031   0.873759039650446   0.02860181540699222   0.8341259141584701   0.3185610680679547   0.5003608063748556   0.6168270457510014   0.4731701937571937   0.011249739034985004   0.0929707224157336   0.6338496383582116   0.6826772094471524   0.6647934239647546   0.003503799301123841   0.5238094275538544   0.6451192103719835   0.29000408104377223   0.8261720826322685   0.33570841939203494   0.6122038934492646   0.714055200946712   0.8785072532404257   0.20614652497153488   0.25879679790511784   0.8554291196046809   0.004748213589979697   0.17754470956454266   0.42467088374664774   0.5368680515367262   0.5043874072151241   0.5607176638135412   0.951500689989454   0.5256183125017413   0.4114166847993905   0.9268680254553295   0.26882348054230165   0.8608248885369867   0.4079128854982666   0.4030585979014751   0.6237042701703182   0.5708208074932144   0.5817408028659982   0.06735017850944014
0.011500376721053564   0.8567656065465025   0.7032335496255724   0.8612036535379053   0.7527035788159357   0.0013364869418214483   0.6984853360355927   0.6836589439733626   0.32803269506928795   0.4644684354050952   0.19409792882046864   0.12294128015982139   0.3765320050798339   0.9388501229033539   0.7826812440210782   0.19607325470449183   0.10770852453753225   0.07802523436636728   0.37476835852281154   0.7930146568030167   0.48400425436721406   0.5072044268731528   0.7930275556568135   0.7256644782935766   0.47250387764616053   0.6504388203266505   0.08979400603124106   0.8644608247556713   0.7198002988302248   0.6491023333848289   0.39130866999564834   0.18080188078230877   0.39176760376093683   0.18463389797973379   0.1972107411751797   0.05786060062248738   0.015235598681102889   0.24578377507637988   0.41452949715410153   0.8617873459179956   0.9075270741435706   0.1677585407100126   0.039761138631289966   0.0687726891149788   0.4235228197763566   0.6605541138368598   0.2467335829744765   0.3431082108214022   0.951018942130196   0.010115293510209322   0.15693957694323546   0.4786473860657308   0.23121864329997124   0.36101296012538037   0.7656309069475871   0.2978455052834221   0.8394510395390344   0.17637906214564655   0.5684201657724074   0.2399849046609347   0.8242154408579315   0.9305952870692666   0.15389066861830586   0.37819755874293914
0.9166883667143609   0.7628367463592541   0.11412952998701589   0.30942486962796034   0.49316554693800435   0.10228263252239433   0.8673959470125394   0.9663166588065581   0.5421466048078083   0.09216733901218502   0.710456370069304   0.48766927274082733   0.310927961507837   0.7311543788868047   0.9448254631217168   0.18982376745740526   0.47147692196880264   0.5547753167411581   0.37640529734930944   0.9498388627964706   0.6472614811108711   0.6241800296718915   0.22251462873100358   0.5716413040535314   0.7305731143965102   0.8613432833126373   0.10838509874398768   0.2622164344255711   0.23740756745850586   0.759060650790243   0.2409891517314483   0.29589977561901293   0.6952609626506976   0.666893311778058   0.5305327816621443   0.8082305028781855   0.3843330011428605   0.9357389328912533   0.5857073185404276   0.6184067354207804   0.9128560791740579   0.3809636161500952   0.2093020211911181   0.6685678726243098   0.2655945980631868   0.7567835864782038   0.9867873924601145   0.09692656857077837   0.5350214836666766   0.8954403031655664   0.8784022937161269   0.8347101341452073   0.29761391620817074   0.1363796523753234   0.6374131419846786   0.5388103585261944   0.6023529535574732   0.4694863405972654   0.10688036032253419   0.7305798556480088   0.21801995241461267   0.533747407706012   0.5211730417821067   0.11217312022722845
0.3051638732405548   0.15278379155591681   0.3118710205909886   0.44360524760291864   0.039569275177368   0.39600020507771305   0.32508362813087405   0.3466786790321403   0.5045477915106914   0.5005599019121466   0.4466813344147472   0.511968544886933   0.20693387530252066   0.3641802495368232   0.8092681924300686   0.9731581863607386   0.6045809217450475   0.8946939089395578   0.7023878321075344   0.24257833071272983   0.38656096933043477   0.36094650123354577   0.18121479032542778   0.13040521048550138   0.08139709608988   0.20816270967762898   0.8693437697344393   0.6867999628825827   0.041827820912512   0.8121625045999159   0.5442601416035652   0.34012128385044244   0.5372800294018206   0.3116026026877693   0.09757880718881799   0.8281527389635094   0.3303461540992999   0.9474223531509461   0.28831061475874936   0.8549945526027708   0.7257652323542525   0.05272844421138827   0.5859227826512149   0.612416221890041   0.3392042630238177   0.6917819429778425   0.4047079923257871   0.4820110114045396   0.2578071669339377   0.4836192333002135   0.5353642225913479   0.7952110485219569   0.21597934602142568   0.6714567287002976   0.9911040809877827   0.4550897646715145   0.678699316619605   0.35985412601252825   0.8935252737989646   0.626937025708005   0.3483531625203051   0.41243177286158217   0.6052146590402153   0.7719424731052342
0.6225879301660527   0.3597033286501939   0.01929187638900046   0.15952625121519323   0.283383667142235   0.6679213856723514   0.6145838840632134   0.6775152398106536   0.02557650020829736   0.1843021523721379   0.07921966147186553   0.8823041912886966   0.8095971541868717   0.5128454236718404   0.08811558048408286   0.4272144266171822   0.1308978375672666   0.15299129765931208   0.19459030668511818   0.8002774009091771   0.7825446750469615   0.7405595247977299   0.5893756476449028   0.028334927803942873   0.15995674488090875   0.380856196147536   0.5700837712559024   0.8688086765887496   0.8765730777386738   0.7129348104751846   0.955499887192689   0.19129343677809604   0.8509965775303764   0.5286326581030467   0.8762802257208234   0.3089892454893994   0.04139942334350468   0.015787234431206384   0.7881646452367406   0.8817748188722172   0.9105015857762381   0.8627959367718943   0.5935743385516224   0.08149741796304005   0.12795691072927662   0.12223641197416439   0.004198690906719594   0.05316249015909718   0.9680001658483679   0.7413802158266284   0.4341149196508172   0.18435381357034755   0.09142708810969415   0.028445405351443732   0.4786150324581282   0.9930603767922515   0.24043051057931777   0.499812747248397   0.6023348067373048   0.6840711313028521   0.19903108723581311   0.48402551281719064   0.8141701615005641   0.8022963124306349
0.288529501459575   0.6212295760452963   0.2205958229489417   0.7207988944675949   0.1605725907302984   0.4989931640711319   0.2163971320422221   0.6676364043084978   0.19257242488193052   0.7576129482445035   0.7822822123914048   0.4832825907381502   0.10114533677223639   0.7291675428930599   0.3036671799332767   0.4902222139458987   0.8607148261929186   0.22935479564466285   0.701332373195972   0.8061510826430466   0.6616837389571055   0.7453292828274722   0.8871622116954078   0.003854770212411566   0.37315423749753046   0.12409970678217588   0.6665663887464661   0.28305587574481667   0.21258164676723207   0.6251065427110439   0.450169256704244   0.6154194714363189   0.020009221885301545   0.8674935944665404   0.6678870443128392   0.13213688069816867   0.9188638851130652   0.13832605157348052   0.3642198643795625   0.6419146667522699   0.058149058920146546   0.9089712559288177   0.6628874911835906   0.8357635841092235   0.396465319963041   0.16364197310134546   0.7757252794881827   0.8319088138968119   0.023311082465510558   0.03954226631916958   0.10915889074171663   0.5488529381519952   0.8107294356982785   0.41443572360812564   0.6589896340374726   0.9334334667156764   0.790720213812977   0.5469421291415852   0.9911025897246335   0.8012965860175076   0.8718563286999118   0.40861607756810475   0.626882725345071   0.15938191926523768
0.8137072697797653   0.4996448216392871   0.9639952341614805   0.32361833515601424   0.4172419498167242   0.3360028485379416   0.18826995467329768   0.49170952125920236   0.39393086735121363   0.29646058221877203   0.07911106393158104   0.9428565831072071   0.5832014316529351   0.8820248586106464   0.42012142989410844   0.009423116391530777   0.7924812178399582   0.33508272946906115   0.429018840169475   0.20812653037402312   0.9206248891400465   0.9264666519009565   0.8021361148244041   0.04874461110878545   0.10691761936028121   0.42682183026166937   0.8381408806629236   0.7251262759527712   0.689675669543557   0.09081898172372774   0.6498709259896259   0.23341675469356887   0.29574480219234334   0.7943583995049557   0.5707598620580449   0.29056017158636177   0.7125433705394082   0.9123335408943093   0.1506384321639364   0.28113705519483095   0.92006215269945   0.5772508114252481   0.7216195919944615   0.07301052482080785   0.9994372635594035   0.6507841595242918   0.9194834771700574   0.024265913712022396   0.8925196441991223   0.22396232926262244   0.08134259650713384   0.2991396377592512   0.2028439746555653   0.1331433475388947   0.43147167051750795   0.06572288306568232   0.9070991724632219   0.338784948033939   0.860711808459463   0.7751627114793206   0.19455580192381375   0.42645140713962965   0.7100733762955267   0.4940256562844896
0.27449364922436376   0.8492005957143814   0.9884537843010652   0.42101513146368175   0.27505638566496027   0.19841643619008967   0.06897030713100784   0.39674921775165933   0.38253674146583794   0.9744541069274673   0.987627710623874   0.09760957999240819   0.17969276681027263   0.8413107593885725   0.5561560401063661   0.03188669692672587   0.27259359434705066   0.5025258113546336   0.6954442316469029   0.2567239854474053   0.07803779242323693   0.07607440421500389   0.9853708553513763   0.7626983291629157   0.8035441431988731   0.22687380850062244   0.996917071050311   0.34168319769923394   0.5284877575339129   0.028457372310532757   0.9279467639193032   0.9449339799475746   0.14595101606807495   0.05400326538306553   0.9403190532954292   0.8473243999551664   0.9662582492578023   0.21269250599449302   0.38416301318906315   0.8154377030284405   0.6936646549107517   0.7101666946398595   0.6887187815421602   0.5587137175810353   0.6156268624875147   0.6340922904248556   0.7033479261907839   0.7960153884181195   0.8120827192886416   0.40721848192423316   0.7064308551404729   0.4543321907188856   0.28359496175472865   0.3787611096137004   0.7784840912211697   0.509398210771311   0.1376439456866537   0.32475784423063486   0.8381650379257405   0.6620738108161446   0.17138569642885138   0.11206533823614186   0.45400202473667733   0.846636107787704
0.4777210415180997   0.4018986435962824   0.7652832431945171   0.2879223902066688   0.8620941790305849   0.7678063531714268   0.06193531700373326   0.4919070017885493   0.05001145974194341   0.36058787124719366   0.35550446186326035   0.03757481106966369   0.7664164979872148   0.9818267616334933   0.5770203706420907   0.5281766002983527   0.6287725523005611   0.6570689174028584   0.7388553327163502   0.8661027894822081   0.4573868558717097   0.5450035791667166   0.28485330797967284   0.019466681694504103   0.97966581435361   0.1431049355704342   0.5195700647851557   0.7315442914878353   0.11757163532302496   0.3752985823990074   0.4576347477814224   0.23963728969928602   0.06756017558108156   0.014710711151813707   0.10213028591816202   0.20206247862962234   0.3011436775938668   0.032883949518320424   0.5251099152760713   0.6738858783312697   0.6723711252933058   0.375815032115462   0.7862545825597211   0.8077830888490615   0.21498426942159612   0.8308114529487455   0.5014012745800484   0.7883164071545574   0.23531845506798615   0.6877065173783112   0.9818312097948927   0.056772115666722085   0.11774681974496119   0.31240793497930386   0.5241964620134704   0.817134825967436   0.05018664416387964   0.29769722382749014   0.4220661760953083   0.6150723473378137   0.7490429665700128   0.26481327430916973   0.896956260819237   0.9411864690065441
0.07667184127670705   0.8889982421937077   0.11070167825951578   0.13340338015748257   0.8616875718551109   0.058186789244962296   0.6093004036794675   0.3450869730029252   0.6263691167871248   0.37048027186665106   0.6274691938845747   0.2883148573362031   0.5086222970421636   0.058072336887347184   0.10327273187110439   0.47118003136876707   0.4584356528782839   0.760375113059857   0.6812065557757961   0.8561076840309534   0.7093926863082711   0.49556183875068727   0.7842502949565592   0.9149212150244093   0.632720845031564   0.6065635965569796   0.6735486166970434   0.7815178348669267   0.7710332731764531   0.5483768073120172   0.06424821301757594   0.4364308618640015   0.14466415638932836   0.1778965354453662   0.4367790191330012   0.14811600452779838   0.6360418593471648   0.11982419855801901   0.33350628726189685   0.6769359731590313   0.17760620646888087   0.359449085498162   0.6522997314861008   0.820828289128078   0.46821352016060974   0.8638872467474747   0.8680494365295416   0.9059070741036688   0.8354926751290457   0.25732365019049513   0.19450081983249823   0.12438923923674207   0.06445940195259259   0.7089468428784779   0.1302526068149223   0.6879583773727406   0.9197952455632642   0.5310503074331117   0.693473587681921   0.5398423728449422   0.28375338621609947   0.4112261088750927   0.3599673004200242   0.8629063996859109
0.10614717974721859   0.05177702337693069   0.7076675689339235   0.042078110557832886   0.6379336595866089   0.187889776629456   0.8396181324043819   0.13617103645416415   0.8024409844575631   0.9305661264389609   0.6451173125718836   0.011781797217422084   0.7379815825049705   0.22161928356048294   0.5148647057569613   0.3238234198446815   0.8181863369417063   0.6905689761273712   0.8213911180750403   0.7839810469997393   0.5344329507256068   0.2793428672522785   0.46142381765501606   0.9210746473138284   0.42828577097838827   0.22756584387534784   0.7537562487210926   0.8789965367559955   0.7903521113917794   0.03967606724589185   0.9141381163167107   0.7428255003018314   0.9879111269342163   0.10910994080693102   0.26902080374482706   0.7310437030844094   0.2499295444292458   0.887490657246448   0.7541560979878658   0.4072202832397278   0.4317432074875395   0.19692168111907687   0.9327649799128255   0.6232392362399886   0.8973102567619327   0.9175788138667983   0.4713411622578094   0.7021645889261601   0.46902448578354444   0.6900129699914505   0.7175849135367168   0.8231680521701645   0.678672374391765   0.6503369027455587   0.8034467972200061   0.08034255186833315   0.6907612474575486   0.5412269619386276   0.534425993475179   0.34929884878392387   0.4408317030283028   0.6537363046921796   0.7802698954873133   0.942078565544196
0.009088495540763273   0.45681462357310265   0.8475049155744879   0.31883932930420755   0.11177823877883059   0.5392358097063044   0.37616375331667845   0.6166747403780475   0.6427537529952861   0.8492228397148538   0.6585788397799616   0.793506688207883   0.9640813786035212   0.19888593696929513   0.8551320425599555   0.7131641363395498   0.2733201311459726   0.6576589750306675   0.32070604908477635   0.3638652875556259   0.8324884281176698   0.003922670338487979   0.540436153597463   0.42178672201142986   0.8233999325769065   0.5471080467653853   0.6929312380229751   0.10294739270722231   0.7116216937980759   0.007872237059081017   0.3167674847062967   0.4862726523291748   0.06886794080278974   0.15864939734422723   0.6581886449263351   0.6927659641212919   0.10478656219926853   0.9597634603749321   0.8030566023663797   0.9796018277817422   0.831466431053296   0.30210448534426454   0.4823505532816033   0.6157365402261162   0.9989780029356262   0.29818181500577656   0.9419143996841403   0.1939498182146864   0.17557807035871972   0.7510737682403913   0.2489831616611652   0.09100242550746408   0.4639563765606438   0.7432015311813103   0.9322156769548685   0.6047297731782892   0.3950884357578541   0.584552133837083   0.2740270320285334   0.9119638090569974   0.29030187355858555   0.624788673462151   0.47097042966215374   0.9323619812752552
0.45883544250528957   0.3226841881178864   0.9886198763805505   0.3166254410491389   0.45985743956966335   0.024502373112109805   0.04670547669641016   0.12267562283445252   0.28427936921094366   0.27342860487171855   0.7977223150352449   0.03167319732698843   0.8203229926502998   0.5302270736904083   0.8655066380803764   0.4269434241486992   0.42523455689244577   0.9456749398533253   0.591479606051843   0.5149796150917019   0.13493268333386024   0.32088626639117435   0.12050917638968929   0.5826176338164467   0.6760972408285707   0.9982020782732879   0.13188930000913882   0.2659921927673078   0.2162398012589073   0.9736997051611781   0.08518382331272867   0.14331656993285527   0.9319604320479636   0.7002711002894596   0.2874615082774837   0.11164337260586683   0.1116374393976638   0.1700440265990513   0.4219548701971072   0.6846999484571676   0.686402882505218   0.224369086745726   0.8304752641452642   0.1697203333654658   0.5514701991713578   0.9034828203545516   0.7099660877555749   0.5871026995490191   0.875372958342787   0.9052807420812637   0.578076787746436   0.3211105067817113   0.6591331570838798   0.9315810369200856   0.49289296443370734   0.17779393684885605   0.7271727250359161   0.23130993663062602   0.20543145615622369   0.06615056424298921   0.6155352856382523   0.06126591003157474   0.7834765859591165   0.38145061578582157
0.9291324031330344   0.8368968232858487   0.9530013218138523   0.21173028242035577   0.3776622039616766   0.9334140029312971   0.24303523405827746   0.6246275828713367   0.5022892456188894   0.028133260850033315   0.6649584463118414   0.30351707608962536   0.8431560885350097   0.0965522239299477   0.17206548187813406   0.1257231392407693   0.11598336349909352   0.8652422872993216   0.9666340257219104   0.059572574997780105   0.5004480778608411   0.803976377267747   0.18315743976279392   0.6781219592119585   0.5713156747278068   0.9670795539818982   0.2301561179489416   0.46639167679160276   0.1936534707661302   0.033665551050601136   0.9871208838906641   0.8417640939202661   0.6913642251472407   0.005532290200567826   0.32216243757882274   0.5382470178306408   0.848208136612231   0.9089800662706201   0.15009695570068865   0.41252387858987144   0.7322247731131375   0.04373777897129845   0.18346292997877825   0.35295130359209137   0.23177669525229636   0.2397614017035515   0.00030549021598433464   0.6748293443801328   0.6604610205244895   0.2726818477216533   0.7701493722670427   0.20843766758853   0.46680754975835936   0.23901629667105218   0.7830284883763786   0.36667357366826386   0.7754433246111186   0.23348400647048434   0.4608660507975558   0.8284265558376231   0.9272351879988876   0.3245039401998642   0.3107690950968672   0.4159026772477517
0.19501041488575005   0.2807661612285658   0.12730616511808893   0.06295137365566034   0.9632337196334537   0.04100475952501427   0.1270006749021046   0.3881220292755275   0.30277269910896415   0.768322911803361   0.3568513026350619   0.17968436168699753   0.8359651493506048   0.5293066151323088   0.5738228142586833   0.8130107880187336   0.060521824739486176   0.2958226086618244   0.11295676346112746   0.9845842321811106   0.1332866367405986   0.9713186684619601   0.8021876683642603   0.5686815549333588   0.9382762218548486   0.6905525072333945   0.6748815032461714   0.5057301812776985   0.9750425022213949   0.6495477477083801   0.5478808283440667   0.11760815200217095   0.6722698031124307   0.8812248359050192   0.19102952570900486   0.9379237903151734   0.836304653761826   0.3519182207727104   0.6172067114503216   0.12491300229643977   0.7757828290223397   0.056095612110886005   0.5042499479891941   0.14032877011532924   0.6424961922817412   0.08477694364892582   0.7020622796249338   0.5716472151819704   0.7042199704268925   0.3942244364155314   0.027180776378762518   0.0659170339042719   0.7291774682054978   0.7446766887071513   0.4792999480346958   0.9483088819021009   0.056907665093067   0.8634518528021321   0.2882704223256909   0.010385091586927521   0.22060301133124108   0.5115336320294217   0.6710637108753693   0.8854720892904877
0.4448201823089013   0.45543801991853566   0.16681376288617525   0.7451433191751585   0.8023239900271601   0.3706610762696098   0.4647514832612414   0.1734961039931881   0.09810401960026757   0.9764366398540785   0.43757070688247884   0.1075790700889162   0.3689265513947698   0.23175995114692716   0.9582707588477831   0.15927018818681526   0.3120188863017028   0.36830809834479505   0.6700003365220921   0.14888509659988775   0.09141587497046177   0.8567744663153735   0.9989366256467228   0.2634130073094   0.6465956926615605   0.40133644639683774   0.8321228627605476   0.5182696881342415   0.8442717026344003   0.030675370127227927   0.3673713794993062   0.34477358414105336   0.7461676830341327   0.054238730273149495   0.9298006726168273   0.23719451405213718   0.3772411316393629   0.8224787791262224   0.9715299137690442   0.0779243258653219   0.06522224533766005   0.45417068078142725   0.30152957724695206   0.9290392292654341   0.9738063703671983   0.5973962144660538   0.30259295160022925   0.6656262219560342   0.32721067770563783   0.19605976806921607   0.47047008883968167   0.14735653382179265   0.4829389750712375   0.16538439794198814   0.10309870934037545   0.8025829496807393   0.7367712920371048   0.11114566766883865   0.17329803672354813   0.5653884356286021   0.3595301603977419   0.2886668885426163   0.2017681229545039   0.4874641097632802
0.29430791506008186   0.834496207761189   0.9002385457075518   0.5584248804978461   0.32050154469288356   0.2370999932951352   0.5976455941073225   0.892798658541812   0.9932908669872458   0.04104022522591913   0.12717550526764093   0.7454421247200193   0.5103518919160083   0.875655827283931   0.024076795927265485   0.94285917503928   0.7735805998789035   0.7645101596150923   0.8507787592037174   0.3774707394106779   0.41405043948116155   0.475843271072476   0.6490106362492135   0.8900066296473976   0.11974252442107972   0.641347063311287   0.7487720905416617   0.3315817491495516   0.7992409797281962   0.40424707001615173   0.1511264964343391   0.4387830906077397   0.8059501127409504   0.36320684479023263   0.02395099116669816   0.6933409658877204   0.2955982208249422   0.48755101750630164   0.9998741952394327   0.7504817908484404   0.5220176209460388   0.7230408578912093   0.14909543603571532   0.37301105143776253   0.10796718146487719   0.2471975868187333   0.5000847997865018   0.48300442179036485   0.9882246570437975   0.6058505235074464   0.7513127092448402   0.15142267264081324   0.1889836773156013   0.2016034534912946   0.6001862128105011   0.7126395820330735   0.38303356457465093   0.838396608701062   0.5762352216438029   0.019298616145353168   0.08743534374970874   0.3508455911947604   0.5763610264043703   0.26881682529691275
0.56541772280367   0.627804733303551   0.4272655903686549   0.8958057738591503   0.4574505413387928   0.3806071464848178   0.9271807905821531   0.4128013520687854   0.46922588429499534   0.7747566229773715   0.17586808133731296   0.26137867942797216   0.280242206979394   0.5731531694860769   0.5756818685268119   0.5487390973948986   0.8972086424047431   0.7347565607850148   0.999446646883009   0.5294404812495455   0.8097732986550343   0.38391096959025445   0.4230856204786388   0.26062365595263265   0.24435557585136436   0.7561062362867034   0.9958200301099839   0.3648178820934824   0.7869050345125715   0.3754990898018856   0.06863923952783077   0.952016530024697   0.3176791502175762   0.6007424668245142   0.8927711581905178   0.6906378505967249   0.037436943238182155   0.02758929733843733   0.3170892896637059   0.1418987532018263   0.14022830083343904   0.2928327365534225   0.3176426427806969   0.6124582719522809   0.3304550021784047   0.9089217669631681   0.8945570223020581   0.3518346159996482   0.08609942632704033   0.15281553067646467   0.8987369921920743   0.9870167339061658   0.2991943918144688   0.7773164408745791   0.8300977526642435   0.03500020388146879   0.9815152415968926   0.17657397405006492   0.9373265944737257   0.3443623532847439   0.9440782983587105   0.1489846767116276   0.6202373048100197   0.20246360008291764
0.8038499975252714   0.8561519401582051   0.30259466202932284   0.5900053281306368   0.4733949953468667   0.947230173195037   0.4080376397272647   0.23817071213098853   0.38729556901982637   0.7944146425185724   0.5093006475351904   0.2511539782248227   0.08810117720535758   0.01709820164399328   0.679202894870947   0.21615377434335395   0.10658593560846497   0.8405242275939283   0.7418763003972213   0.8717914210586101   0.1625076372497545   0.6915395508823008   0.12163899558720158   0.6693278209756924   0.3586576397244831   0.8353876107240956   0.8190443335578788   0.07932249284505563   0.8852626443776164   0.8881574375290586   0.41100669383061406   0.841151780714067   0.49796707535779   0.09374279501048625   0.9017060462954236   0.5899978024892444   0.4098658981524324   0.07664459336649297   0.2225031514244767   0.3738440281458904   0.30327996254396744   0.23612036577256462   0.4806268510272554   0.5020526070872804   0.14077232529421294   0.5445808148902639   0.3589878554400538   0.8327247861115881   0.7821146855697299   0.7091932041661682   0.539943521882175   0.7534022932665324   0.8968520411921135   0.8210357666371095   0.12893682805156093   0.9122505125524653   0.3988849658343234   0.7272929716266233   0.22723078175613728   0.3222527100632209   0.989019067681891   0.6506483782601303   0.00472763033166061   0.9484086819173305
0.6857391051379236   0.4145280124875657   0.5241007793044052   0.4463560748300501   0.5449667798437106   0.8699471975973019   0.16511292386435147   0.6136312887184621   0.7628520942739807   0.16075399343113367   0.6251694019821765   0.8602289954519297   0.8660000530818673   0.3397182267940241   0.49623257393061554   0.9479784828994644   0.4671150872475439   0.6124252551674008   0.2690017921744783   0.6257257728362435   0.47809601956565295   0.9617768769072704   0.26427416184281766   0.677317090918913   0.7923569144277294   0.5472488644197047   0.7401733825384124   0.2309610160888629   0.24739013458401882   0.6773016668224029   0.575060458674061   0.6173297273704008   0.48453804031003805   0.5165476733912692   0.9498910566918845   0.7571007319184712   0.6185379872281708   0.17682944659724512   0.4536584827612689   0.8091222490190068   0.1514228999806268   0.5644041914298443   0.18465669058679066   0.18339647618276322   0.6733268804149739   0.6026273145225739   0.920382528743973   0.5060793852638502   0.8809699659872444   0.05537845010286922   0.1802091462055606   0.27511836917498733   0.6335798314032256   0.37807678328046634   0.6051486875314996   0.6577886418045865   0.14904179109318758   0.8615291098891972   0.6552576308396152   0.9006879098861154   0.5305038038650168   0.6846996632919521   0.2015991480783463   0.09156566086710867
0.37908090388439003   0.12029547186210769   0.016942457491555655   0.9081691846843455   0.7057540234694162   0.5176681573395338   0.09655992874758265   0.4020897994204952   0.8247840574821717   0.4622897072366645   0.9163507825420221   0.1269714302455079   0.19120422607894605   0.08421292395619817   0.3112020950105224   0.4691827884409214   0.04216243498575848   0.222683814067001   0.6559444641709071   0.568494878554806   0.5116586311207416   0.5379841507750489   0.45434531609256085   0.4769292176876973   0.13257772723635158   0.41768867891294126   0.4374028586010052   0.5687600330033519   0.42682370376693546   0.9000205215734075   0.3408429298534225   0.16667023358285665   0.6020396462847637   0.43773081433674293   0.4244921473114005   0.03969880333734878   0.4108354202058177   0.3535178903805448   0.11329005230087813   0.5705160148964274   0.3686729852200592   0.1308340763135438   0.457345588129971   0.0020211363416214093   0.8570143540993176   0.5928499255384948   0.0030002720374101596   0.5250919186539241   0.724436626862966   0.17516124662555357   0.565597413436405   0.9563318856505723   0.29761292309603055   0.2751407250521461   0.22475448358298247   0.7896616520677155   0.6955732768112668   0.8374099107154032   0.8002623362715819   0.7499628487303668   0.2847378566054491   0.48389202033485834   0.6869722839707039   0.17944683383393936
0.91606487138539   0.3530579440213145   0.22962669584073286   0.17742569749231796   0.05905051728607233   0.7602080184828197   0.2266264238033227   0.6523337788383938   0.33461389042310635   0.5850467718572662   0.6610290103669177   0.6960018931878217   0.03700096732707581   0.30990604680512   0.43627452678393525   0.9063402411201061   0.341427690515809   0.4724961360897169   0.6360121905123532   0.15637739238973933   0.056689833910359894   0.9886041157548586   0.9490399065416494   0.9769305585557999   0.14062496252496998   0.635546171733544   0.7194132107009166   0.799504861063482   0.08157444523889765   0.8753381532507244   0.49278678689759386   0.14717108222508812   0.7469605548157913   0.2902913813934582   0.8317577765306762   0.45116918903726644   0.7099595874887155   0.9803853345883382   0.3954832497467409   0.5448289479171603   0.3685318969729065   0.5078891984986212   0.7594710592343876   0.388451555527421   0.3118420630625466   0.5192850827437627   0.8104311526927381   0.41152099697162103   0.1712171005375766   0.8837389110102186   0.0910179419918216   0.6120161359081391   0.08964265529867896   0.008400757759494292   0.5982311550942278   0.4648450536830509   0.34268210048288766   0.7181093763660361   0.7664733785635516   0.013675864645784474   0.6327225129941721   0.7377240417776979   0.37099012881681076   0.4688469167286241
0.2641906160212657   0.2298348432790766   0.6115190695824232   0.08039536120120312   0.9523485529587191   0.7105497605353139   0.801087916889685   0.6688743642295821   0.7811314524211425   0.8268108495250953   0.7100699748978634   0.056858228321443036   0.6914887971224636   0.818410091765601   0.11183881980363561   0.5920131746383921   0.34880669663957586   0.10030071539956491   0.345365441240084   0.5783373099926077   0.7160841836454037   0.362576673621867   0.9743753124232732   0.10949039326398351   0.451893567624138   0.13274183034279044   0.3628562428408501   0.029095032062780374   0.4995450146654189   0.42219206980747653   0.5617683259511651   0.3602206678331983   0.7184135622442764   0.5953812202823813   0.8516983510533018   0.30336243951175523   0.026924765121812886   0.7769711285167803   0.7398595312496662   0.7113492648733631   0.678118068482237   0.6766704131172154   0.3944940900095822   0.1330119548807555   0.9620338848368333   0.31409373949534836   0.4201187775863089   0.02352156161677201   0.5101403172126953   0.1813519091525579   0.05726253474545879   0.9944265295539917   0.010595302547276395   0.7591598393450814   0.4954942087942936   0.6342058617207933   0.292181740303   0.16377861906270008   0.6437958577409918   0.3308434222090381   0.26525697518118707   0.3868074905459198   0.9039363264913257   0.6194941573356749
0.5871389066989501   0.7101370774287044   0.5094422364817435   0.4864822024549194   0.6251050218621168   0.39604333793335605   0.08932345889543458   0.4629606408381474   0.11496470464942145   0.21469142878079817   0.0320609241499758   0.4685341112841558   0.10436940210214506   0.4555315894357168   0.5365667153556821   0.8343282495633625   0.812187661799145   0.29175297037301673   0.8927708576146903   0.5034848273543243   0.546930686617958   0.9049454798270969   0.9888345311233646   0.8839906700186494   0.9597917799190079   0.19480840239839253   0.47939229464162114   0.39750846756373   0.3346867580568912   0.7987650644650365   0.39006883574618656   0.9345478267255826   0.21972205340746973   0.5840736356842383   0.35800791159621076   0.4660137154414268   0.11535265130532465   0.12854204624852147   0.8214411962405286   0.6316854658780643   0.3031649895061796   0.8367890758755048   0.9286703386258383   0.12820063852373995   0.7562343028882216   0.9318435960484078   0.9398358075024736   0.24420996850509055   0.7964425229692137   0.7370351936500152   0.46044351286085244   0.8467015009413605   0.4617557649123225   0.9382701291849788   0.0703746771146659   0.912153674215778   0.24203371150485278   0.3541964935007405   0.7123667655184551   0.44613995877435125   0.12668106019952813   0.22565444725221903   0.8909255692779265   0.814454492896287
0.8235160706933485   0.3888653713767143   0.9622552306520883   0.686253854372547   0.06728176780512697   0.4570217753283065   0.022419423149614648   0.44204388586745647   0.2708392448359133   0.7199865816782912   0.5619759102887621   0.5953423849260959   0.8090834799235909   0.7817164524933125   0.49160123317409626   0.6831887107103178   0.5670497684187381   0.427519958992572   0.7792344676556412   0.2370487519359666   0.4403687082192099   0.20186551174035294   0.8883088983777147   0.4225942590396796   0.6168526375258614   0.8130001403636387   0.9260536677256264   0.7363404046671326   0.5495708697207344   0.3559783650353322   0.9036342445760117   0.29429651879967617   0.27873162488482106   0.6359917833570409   0.3416583342872495   0.6989541338735803   0.46964814496123025   0.8542753308637284   0.8500571011131532   0.01576542316326237   0.9025983765424922   0.4267553718711565   0.0708226334575121   0.7787166712272957   0.4622296683232823   0.22488986013080353   0.18251373507979748   0.3561224121876161   0.8453770307974209   0.4118897197671649   0.25646006735417115   0.6197820075204835   0.29580616107668645   0.05591135473183269   0.35282582277815944   0.32548548872080735   0.017074536191865355   0.41991957137479174   0.011167488490909946   0.6265313548472271   0.5474263912306351   0.5656442405110633   0.1611103873777567   0.6107659316839648
0.6448280146881429   0.1388888686399068   0.09028775392024463   0.8320492604566689   0.18259834636486066   0.9139990085091033   0.9077740188404472   0.47592684826905285   0.33722131556743984   0.5021092887419384   0.651313951486276   0.8561448407485693   0.04141515449075337   0.4461979340101057   0.29848812870811653   0.530659352027762   0.02434061829888802   0.02627836263531397   0.2873206402172066   0.9041279971805349   0.4769142270682529   0.4606341221242507   0.1262102528394499   0.29336206549657023   0.83208621238011   0.32174525348434385   0.03592249891920525   0.4613128050399013   0.6494878660152493   0.4077462449752406   0.12814848007875812   0.9853859567708485   0.3122665504478095   0.9056369562333022   0.4768345285924821   0.1292411160222791   0.27085139595705615   0.45943902222319644   0.17834639988436557   0.5985817639945171   0.24651077765816812   0.43316065958788247   0.891025759667159   0.6944537668139822   0.7695965505899152   0.9725265374636318   0.764815506827709   0.4010917013174119   0.9375103382098052   0.6507812839792879   0.7288930079085039   0.9397788962775105   0.2880224721945559   0.24303503900404735   0.6007445278297457   0.9543929395066622   0.9757559217467464   0.3373980827707452   0.12390999923726362   0.825151823484383   0.7049045257896902   0.8779590605475487   0.945563599352898   0.2265700594898659
0.4583937481315221   0.4447984009596662   0.054537839685739074   0.5321162926758838   0.688797197541607   0.4722718634960344   0.28972233285802995   0.1310245913584719   0.7512868593318017   0.8214905795167464   0.5608293249495261   0.19124569508096131   0.4632643871372458   0.5784555405126991   0.9600847971197805   0.2368527555742992   0.48750846539049947   0.24105745774195395   0.8361747978825168   0.4117009320899162   0.7826039396008092   0.36309839719440523   0.8906111985296188   0.18513087260005032   0.3242101914692871   0.918299996234739   0.8360733588438797   0.6530145799241666   0.6354129939276801   0.4460281327387046   0.5463510259858497   0.5219899885656947   0.8841261345958784   0.6245375532219581   0.9855217010363235   0.3307442934847334   0.4208617474586326   0.04608201270925907   0.025436903916543147   0.09389153791043417   0.9333532820681332   0.8050245549673051   0.18926210603402635   0.6821906058205179   0.1507493424673239   0.44192615777289984   0.2986509075044076   0.49705973322046765   0.8265391509980368   0.5236261615381608   0.4625775486605279   0.8440451532963011   0.19112615707035666   0.07759802879945617   0.9162265226746782   0.3220551647306064   0.3070000224744782   0.453060475577498   0.9307048216383547   0.991310871245873   0.8861382750158456   0.4069784628682389   0.9052679177218115   0.8974193333354389
0.9527849929477126   0.6019539079009338   0.7160058116877852   0.21522872751492092   0.8020356504803886   0.16002775012803397   0.41735490418337756   0.7181689942944532   0.9754964994823518   0.6364015885898732   0.9547773555228496   0.8741238409981522   0.7843703424119951   0.558803559790417   0.038550832848171415   0.5520686762675457   0.4773703199375169   0.105743084212919   0.10784601120981675   0.5607578050216727   0.5912320449216713   0.6987646213446801   0.20257809348800523   0.6633384716862338   0.6384470519739587   0.09681071344374627   0.48657228180022005   0.44810974417131283   0.8364114014935701   0.9367829633157123   0.06921737761684252   0.7299407498768595   0.8609149020112182   0.30038137472583915   0.11444002209399289   0.8558169088787074   0.07654455959922307   0.7415778149354222   0.07588918924582147   0.30374823261116163   0.5991742396617061   0.6358347307225032   0.9680431780360047   0.742990427589489   0.007942194740034915   0.9370701093778231   0.7654650845479994   0.07965195590325518   0.3694951427660762   0.8402593959340768   0.2788928027477794   0.6315422117319424   0.5330837412725061   0.9034764326183645   0.2096754251309369   0.9016014618550827   0.6721688392612879   0.6030950578925254   0.09523540303694401   0.04578455297637535   0.5956242796620649   0.8615172429571032   0.019346213791122537   0.7420363203652137
0.9964500400003586   0.2256825122346   0.05130303575511781   0.9990458927757248   0.9885078452603238   0.2886124028567769   0.2858379512071183   0.9193939368724695   0.6190127024942476   0.4483530069227001   0.0069451484593389175   0.2878517251405272   0.0859289612217414   0.5448765743043356   0.7972697233284021   0.3862502632854445   0.4137601219604535   0.9417815164118102   0.7020343202914581   0.34046571030906914   0.8181358422983886   0.08026427345470705   0.6826881065003355   0.5984293899438554   0.8216858022980299   0.8545817612201071   0.6313850707452177   0.5993834971681307   0.8331779570377061   0.5659693583633302   0.34554711953809936   0.6799895602956612   0.21416525454345858   0.11761635144063005   0.33860197107876044   0.3921378351551339   0.12823629332171718   0.5727397771362944   0.5413322477503584   0.005887571869689437   0.7144761713612637   0.6309582607244842   0.8392979274589004   0.6654218615606203   0.8963403290628751   0.5506939872697773   0.1566098209585649   0.06699247161676487   0.07465452676484516   0.6961122260496702   0.5252247502133472   0.46760897444863414   0.241476569727139   0.13014286768634004   0.1796776306752479   0.787619414152973   0.027311315183680407   0.01252651624570999   0.8410756595964874   0.3954815789978391   0.8990750218619632   0.4397867391094155   0.29974341184612907   0.3895940071281497
0.1845988505006995   0.8088284783849312   0.46044548438722865   0.7241721455675294   0.28825852143782443   0.258134491115154   0.3038356634286638   0.6571796739507645   0.21360399467297925   0.5620222650654839   0.7786109132153166   0.18957069950213032   0.9721274249458403   0.4318793973791438   0.5989332825400687   0.4019512853491573   0.9448161097621598   0.41935288113343383   0.7578576229435813   0.006469706351318213   0.04574108790019663   0.9795661420240184   0.45811421109745215   0.6168756992231685   0.8611422373994971   0.17073766363908707   0.9976687267102234   0.8927035536556392   0.5728837159616728   0.912603172523933   0.6938330632815597   0.2355238797048747   0.35927972128869345   0.35058090745844916   0.9152221500662432   0.0459531802027444   0.3871522963428532   0.9187015100793053   0.31628886752617447   0.644001894853587   0.44233618658069335   0.49934862894587145   0.5584312445825932   0.6375321885022689   0.39659509868049675   0.5197824869218531   0.10031703348514108   0.020656489279100323   0.5354528612809996   0.3490448232827661   0.10264830677491758   0.1279529356234611   0.9625691453193269   0.43644165075883307   0.4088152434933579   0.8924290559185863   0.6032894240306335   0.0858607433003839   0.4935930934271147   0.846475875715842   0.21613712768778023   0.1671592332210786   0.17730422590094028   0.2024739808622549
0.7738009411070869   0.6678106042752071   0.618872981318347   0.564941792359986   0.3772058424265901   0.14802811735335394   0.5185559478332059   0.5442853030808857   0.8417529811455905   0.7989832940705879   0.41590764105828837   0.4163323674574246   0.8791838358262637   0.3625416433117548   0.007092397564930486   0.5239033115388382   0.27589441179563023   0.2766809000113709   0.5134993041378157   0.6774274358229961   0.059757284107849994   0.10952166679029232   0.3361950782368755   0.47495345496074126   0.2859563430007631   0.44171106251508524   0.7173220969185284   0.9100116626007553   0.908750500574173   0.29368294516173127   0.19876614908532247   0.36572635951986954   0.06699751942858245   0.4946996510911434   0.7828585080270342   0.949393992062445   0.18781368360231881   0.1321580077793886   0.7757661104621036   0.4254906805236068   0.9119192718066886   0.8554771077680177   0.2622668063242879   0.7480632447006106   0.8521619876988386   0.7459554409777254   0.9260717280874124   0.2731097897398693   0.5662056446980754   0.30424437846264013   0.20874963116888395   0.36309812713911405   0.6574551441239025   0.01056143330090887   0.009983482083561484   0.9973717676192445   0.59045762469532   0.5158617822097654   0.22712497405652737   0.04797777555679954   0.4026439410930012   0.38370377443037684   0.45135886359442373   0.6224870950331928
0.49072466928631264   0.5282266666623592   0.18909205727013587   0.8744238503325822   0.638562681587474   0.7822712256846338   0.26302032918272344   0.6013140605927129   0.07235703688939855   0.4780268472219937   0.05427069801383949   0.23821593345359882   0.41490189276549605   0.4674654139210848   0.044287215930278005   0.2408441658343543   0.824444268070176   0.9516036317113193   0.8171622418737506   0.19286639027755478   0.42180032697717484   0.5678998572809425   0.3658033782793269   0.570379295244362   0.9310756576908622   0.03967319061858329   0.176711321009191   0.6959554449117799   0.29251297610338817   0.25740196493394946   0.9136909918264675   0.09464138431906696   0.22015593921398963   0.7793751177119558   0.8594202938126281   0.8564254508654682   0.8052540464484935   0.311909703790871   0.8151330778823501   0.6155812850311139   0.9808097783783175   0.3603060720795517   0.9979708360085995   0.42271489475355906   0.5590094514011427   0.7924062147986092   0.6321674577292725   0.852335599509197   0.6279337937102805   0.752733024180026   0.4554561367200815   0.1563801545974172   0.3354208176068923   0.49533105924607645   0.5417651448936139   0.06173877027835023   0.11526487839290268   0.7159559415341207   0.6823448510809859   0.20531331941288208   0.31001083194440915   0.4040462377432496   0.8672117731986358   0.5897320343817682
0.32920105356609164   0.04374016566369792   0.8692409371900364   0.16701713962820922   0.770191602164949   0.2513339508650887   0.23707347946076382   0.31468154011901217   0.14225780845466846   0.4986009266850628   0.7816173427406823   0.15830138552159498   0.8068369908477762   0.003269867438986303   0.23985219784706835   0.09656261524324476   0.6915721124548735   0.28731392590486565   0.5575073467660825   0.8912492958303627   0.38156128051046434   0.883267688161616   0.6902955735674466   0.3015172614485944   0.052360226944372736   0.8395275224979182   0.8210546363774103   0.1345001218203852   0.2821686247794238   0.5881935716328295   0.5839811569166464   0.819818581701373   0.13991081632475533   0.08959264494776667   0.8023638141759641   0.661517196179778   0.33307382547697917   0.08632277750878037   0.5625116163288958   0.5649545809365333   0.6415017130221057   0.7990088516039147   0.005004269562813338   0.6737052851061706   0.25994043251164134   0.9157411634422986   0.31470869599536666   0.3721880236575762   0.20758020556726858   0.07621364094438053   0.4936540596179564   0.237687901837191   0.9254115807878448   0.4880200693115511   0.90967290270131   0.41786932013581796   0.7855007644630895   0.3984274243637844   0.10730908852534574   0.7563521239560399   0.4524269389861103   0.31210464685500405   0.5447974721964499   0.19139754301950665
0.8109252259640046   0.5130957952510894   0.5397932026336366   0.5176922579133361   0.5509847934523633   0.5973546318087907   0.22508450663826993   0.14550423425575987   0.3434045878850947   0.5211409908644101   0.7314304470203136   0.9078163324185688   0.4179930070972499   0.03312092155285908   0.8217575443190036   0.4899470122827509   0.6324922426341604   0.6346934971890746   0.7144484557936579   0.733594888326711   0.18006530364805012   0.3225888503340706   0.16965098359720795   0.5421973453072043   0.36914007768404555   0.8094930550829812   0.6298577809635714   0.024505087393868294   0.8181552842316823   0.21213842327419052   0.40477327432530147   0.8790008531381084   0.47475069634658756   0.6909974324097804   0.673342827304988   0.9711845207195395   0.056757689249337696   0.6578765108569212   0.8515852829859842   0.48123750843678864   0.4242654466151773   0.02318301366784661   0.1371368271923264   0.7476426201100776   0.24420014296712714   0.700594163333776   0.9674858435951185   0.2054452748028733   0.8750600652830816   0.8911011082507948   0.33762806263154704   0.180940187409005   0.05690478105139935   0.6789626849766043   0.9328547883062456   0.3019393342708966   0.5821540847048118   0.9879652525668239   0.2595119610012577   0.330754813551357   0.5253963954554741   0.33008874170990266   0.4079266780152734   0.8495173051145684
0.1011309488402968   0.30690572804205607   0.27078985082294704   0.10187468500449075   0.8569308058731697   0.6063115647082801   0.3033040072278286   0.8964294102016175   0.981870740590088   0.7152104564574853   0.9656759445962816   0.7154892227926125   0.9249659595386888   0.03624777148088097   0.03282115629003597   0.41354988852171587   0.34281187483387693   0.04828251891405705   0.7733091952887783   0.08279507497035887   0.8174154793784029   0.7181937772041543   0.3653825172735049   0.2332777698557905   0.716284530538106   0.4112880491620983   0.09459266645055789   0.13140308485129973   0.8593537246649364   0.8049764844538183   0.7912886592227293   0.23497367464968227   0.8774829840748484   0.08976602799633307   0.8256127146264477   0.5194844518570698   0.9525170245361596   0.053518256515452105   0.7927915583364118   0.10593456333535392   0.6097051497022826   0.005235737601395058   0.019482363047633445   0.023139488364995048   0.7922896703238798   0.28704196039724067   0.6540998457741285   0.7898617185092046   0.07600513978577375   0.8757539112351423   0.5595071793235706   0.6584586336579048   0.21665141512083735   0.07077742678132402   0.7682185201008414   0.4234849590082226   0.33916843104598904   0.981011398784991   0.9426058054743937   0.9040005071511528   0.38665140650982943   0.9274931422695388   0.14981424713798192   0.7980659438157989
0.7769462568075467   0.9222574046681438   0.1303318840903485   0.7749264554508039   0.9846565864836669   0.6352154442709032   0.4762320383162199   0.9850647369415992   0.9086514466978932   0.7594615330357608   0.9167248589926492   0.3266061032836944   0.6920000315770558   0.6886841062544368   0.1485063388918079   0.9031211442754719   0.35283160053106677   0.7076727074694458   0.2059005334174142   0.9991206371243191   0.9661801940212373   0.7801795651999069   0.056086286279432296   0.2010546933085202   0.1892339372136906   0.8579221605317632   0.9257544021890838   0.42612823785771636   0.20457735073002367   0.22270671626086003   0.4495223638728639   0.4410635009161171   0.2959259040321305   0.4632451832250992   0.5327975048802146   0.11445739763242276   0.6039258724550747   0.7745610769706625   0.38429116598840674   0.21133625335695094   0.25109427192400785   0.06688836950121668   0.17839063257099252   0.21221561623263188   0.28491407790277046   0.28670880430130974   0.12230434629156021   0.0111609229241117   0.09568014068907986   0.42878664376954656   0.1965499441024764   0.5850326850663953   0.8911027899590562   0.20607992750868656   0.7470275802296125   0.14396918415027815   0.5951768859269257   0.7428347442835873   0.2142300753493979   0.029511786517855403   0.9912510134718511   0.9682736673129249   0.8299389093609911   0.8181755331609044
0.7401567415478432   0.9013852978117081   0.6515482767899986   0.6059599169282726   0.4552426636450727   0.6146764935103983   0.5292439304984384   0.5947989940041609   0.35956252295599284   0.1858898497408518   0.33269398639596204   0.009766308937765554   0.46845973299693666   0.9798099222321652   0.5856664061663496   0.8657971247874874   0.873282847070011   0.23697517794857795   0.37143633081695165   0.836285338269632   0.88203183359816   0.2687015106356531   0.5414974214559605   0.01810980510872753   0.14187509205031673   0.367316212823945   0.8899491446659619   0.41214988818045495   0.686632428405244   0.7526397193135467   0.36070521416752344   0.8173508941762941   0.32706990544925113   0.5667498695726948   0.028011227771561405   0.8075845852385285   0.8586101724523145   0.5869399473405296   0.4423448216052119   0.9417874604510411   0.9853273253823035   0.34996476939195165   0.07090849078826025   0.10550212218140916   0.10329549178414357   0.08126325875629851   0.5294110693322998   0.08739231707268162   0.9614203997338269   0.7139470459323535   0.6394619246663379   0.6752424288922266   0.27478797132858285   0.9613073266188068   0.2787567104988145   0.8578915347159326   0.9477180658793317   0.394557457046112   0.2507454827272531   0.05030694947740403   0.08910789342701722   0.8076175097055824   0.8084006611220412   0.10851948902636288
0.10378056804471372   0.45765274031363073   0.737492170333781   0.0030173668449537273   0.0004850762605701515   0.3763894815573322   0.2080811010014812   0.9156250497722721   0.03906467652674331   0.6624424356249787   0.5686191763351433   0.24038262088004544   0.7642767051981605   0.7011351090061719   0.28986246583632874   0.38249108616411287   0.8165586393188288   0.3065776519600599   0.03911698310907568   0.3321841366867088   0.7274507458918116   0.4989601422544775   0.23071632198703448   0.22366464766034594   0.6236701778470979   0.04130740194084678   0.4932241516532535   0.22064728081539223   0.6231851015865277   0.6649179203835146   0.2851430506517723   0.3050222310431201   0.5841204250597843   0.00247548475853582   0.7165238743166291   0.06463961016307469   0.819843719861624   0.30134037575236394   0.4266614084803003   0.6821485239989619   0.0032850805427951336   0.994762723792304   0.38754442537122463   0.349964387312253   0.27583433465098356   0.4958025815378265   0.15682810338419015   0.12629973965190705   0.6521641568038857   0.4544951795969797   0.6636039517309367   0.9056524588365148   0.028979055217358052   0.7895772592134651   0.3784609010791643   0.6006302277933947   0.44485863015757365   0.7871017744549293   0.6619370267625352   0.5359906176303201   0.6250149102959498   0.4857613987025654   0.23527561828223492   0.8538420936313582
0.6217298297531546   0.4909986749102614   0.8477311929110103   0.5038777063191052   0.34589549510217105   0.9951960933724349   0.6909030895268201   0.3775779666671982   0.6937313382982854   0.5407009137754551   0.027299137795883527   0.4719255078306833   0.6647522830809273   0.75112365456199   0.6488382367167193   0.8712952800372886   0.21989365292335358   0.9640218801070607   0.986901209954184   0.33530466240696855   0.5948787426274038   0.47826048140449523   0.7516255916719491   0.4814625687756104   0.9731489128742492   0.9872618064942339   0.9038943987609388   0.9775848624565051   0.6272534177720781   0.9920657131217989   0.21299130923411858   0.600006895789307   0.9335220794737928   0.45136479934634377   0.18569217143823508   0.1280813879586237   0.2687697963928656   0.7002411447843537   0.5368539347215159   0.2567861079213351   0.04887614346951197   0.736219264677293   0.5499527247673318   0.9214814455143665   0.45399740084210816   0.25795878327279786   0.7983271330953828   0.44001887673875617   0.48084848796785895   0.270696976778564   0.894432734334444   0.462434014282251   0.8535950701957808   0.27863126365676505   0.6814414251003255   0.862427118492944   0.920072990721988   0.8272664643104213   0.4957492536620904   0.7343457305343203   0.6513031943291224   0.12702531952606752   0.9588953189405746   0.4775596226129852
0.6024270508596105   0.39080605484877445   0.4089425941732427   0.5560781770986187   0.1484296500175023   0.1328472715759766   0.6106154610778599   0.11605930035986255   0.6675811620496434   0.8621502947974126   0.7161827267434159   0.6536252860776116   0.8139860918538625   0.5835190311406475   0.03474130164309043   0.7911981675846675   0.8939131011318746   0.7562525668302262   0.5389920479810001   0.0568524370503473   0.24260990680275213   0.6292272473041587   0.5800967290404255   0.5792928144373621   0.6401828559431417   0.2384211924553843   0.17115413486718278   0.023214637338743405   0.49175320592563937   0.10557392087940769   0.5605386737893229   0.9071553369788808   0.824172043875996   0.24342362608199508   0.844355947045907   0.2535300509012693   0.01018595202213346   0.6599045949413476   0.8096146454028166   0.4623318833166017   0.11627285089025889   0.9036520281111213   0.27062259742181655   0.4054794462662544   0.8736629440875068   0.2744247808069626   0.6905258683813911   0.8261866318288923   0.23348008814436505   0.036003588351578304   0.5193717335142083   0.8029719944901489   0.7417268822187257   0.9304296674721706   0.9588330597248854   0.895816657511268   0.9175548383427297   0.6870060413901755   0.11447711267897837   0.6422866066099987   0.9073688863205962   0.02710144644882798   0.3048624672761618   0.17995472329339704
0.7910960354303374   0.12344941833770667   0.03423986985434527   0.7744752770271427   0.9174330913428306   0.8490246375307441   0.3437140014729542   0.9482886451982504   0.6839530031984655   0.8130210491791658   0.824342267958746   0.14531665070810149   0.9422261209797398   0.8825913817069951   0.8655092082338606   0.24949999319683347   0.02467128263701015   0.19558534031681965   0.7510320955548823   0.6072133865868348   0.11730239631641394   0.16848389386799165   0.4461696282787205   0.42725866329343765   0.32620636088607663   0.04503447553028498   0.4119297584243752   0.6527833862662951   0.40877326954324605   0.1960098379995409   0.06821575695142096   0.7044947410680447   0.7248202663447805   0.38298878882037507   0.24387348899267497   0.5591780903599431   0.7825941453650407   0.5003974071133799   0.37836428075881434   0.30967809716310973   0.7579228627280306   0.3048120667965603   0.6273321852039321   0.702464710576275   0.6406204664116166   0.13632817292856864   0.18116255692521163   0.2752060472828373   0.31441410552554   0.09129369739828365   0.7692327985008365   0.6224226610165423   0.905640835982294   0.8952838593987428   0.7010170415494155   0.9179279199484977   0.18082056963751345   0.5122950705783677   0.4571435525567405   0.3587498295885545   0.39822642427247273   0.011897663464987737   0.07877927179792614   0.04907173242544479
0.6403035615444422   0.7070855966684274   0.4514470865939941   0.3466070218491698   0.9996830951328256   0.5707574237398588   0.2702845296687824   0.07140097456633247   0.6852689896072856   0.4794637263415752   0.501051731167946   0.4489783135497902   0.7796281536249916   0.5841798669428324   0.8000346896185305   0.5310503936012925   0.5988075839874781   0.07188479636446475   0.34289113706179003   0.17230056401273802   0.20058115971500542   0.05998713289947702   0.2641118652638639   0.12322883158729322   0.5602775981705632   0.3529015362310496   0.8126647786698699   0.7766218097381234   0.5605945030377376   0.7821441124911908   0.5423802490010874   0.7052208351717909   0.8753255134304521   0.30268038614961557   0.04132851783314142   0.2562425216220008   0.09569735980546044   0.7185005192067832   0.2412938282146109   0.7251921280207083   0.49688977581798227   0.6466157228423184   0.8984026911528209   0.5528915640079702   0.2963086161029768   0.5866285899428414   0.6342908258889569   0.42966273242067704   0.7360310179324137   0.2337270537117918   0.821626047219087   0.6530409226825536   0.17543651489467596   0.45158294122060105   0.27924579821799966   0.9478200875107626   0.3001110014642239   0.1489025550709855   0.23791728038485824   0.6915775658887618   0.20441364165876347   0.43040203586420234   0.9966234521702474   0.9663854378680536
0.7075238658407812   0.783786313021884   0.09822076101742652   0.41349387386008335   0.4112152497378044   0.19715772307904256   0.4639299351284696   0.9838311414394063   0.6751842318053908   0.9634306693672507   0.6423038879093825   0.3307902187568527   0.4997477169107148   0.5118477281466497   0.3630580896913828   0.38297013124609003   0.1996367154464909   0.3629451730756642   0.12514080930652458   0.6913925653573282   0.9952230737877275   0.9325431372114619   0.1285173571362772   0.7250071274892745   0.2876992079469462   0.14875682418957792   0.030296596118850685   0.31151325362919113   0.8764839582091418   0.9515991011105354   0.5663666609903811   0.3276821121897848   0.20129972640375107   0.9881684317432846   0.9240627730809986   0.9968918934329322   0.7015520094930363   0.4763207035966349   0.5610046833896158   0.6139217621868421   0.5019152940465453   0.11337553052097069   0.43586387408309124   0.922529196829514   0.506692220258818   0.18083239330950882   0.30734651694681403   0.19752206934023944   0.21899301231187177   0.0320755691199309   0.27704992082796337   0.8860088157110483   0.3425090541027299   0.08047646800939554   0.7106832598375823   0.5583267035212635   0.14120932769897887   0.09230803626611095   0.7866204867565836   0.5614348100883314   0.4396573182059426   0.615987332669476   0.22561580336696782   0.9475130479014893
0.9377420241593972   0.5026118021485053   0.7897519292838766   0.024983851071975337   0.43104980390057923   0.32177940883899653   0.4824054123370626   0.8274617817317359   0.21205679158870747   0.28970383971906566   0.2053554915090992   0.9414529660206876   0.8695477374859775   0.2092273717096701   0.49467223167151697   0.38312626249942405   0.7283384097869986   0.11691933544355915   0.7080517449149334   0.8216914524110926   0.28868109158105604   0.5009320027740831   0.4824359415479655   0.8741784045096034   0.35093906742165887   0.9983202006255778   0.6926840122640889   0.8491945534376281   0.9198892635210796   0.6765407917865812   0.21027859992702636   0.02173277170589218   0.7078324719323722   0.38683695206751556   0.004923108417927154   0.08027980568520461   0.8382847344463946   0.1776095803578455   0.5102508767464102   0.6971535431857805   0.109946324659396   0.06069024491428634   0.8021991318314768   0.8754620907746878   0.82126523307834   0.5597582421402032   0.31976319028351136   0.001283686265084456   0.4703261656566811   0.5614380415146255   0.6270791780194225   0.1520891328274564   0.5504369021356015   0.8848972497280443   0.41680057809239607   0.1303563611215642   0.8426044302032293   0.4980602976605287   0.4118774696744689   0.0500765554363596   0.004319695756834663   0.32045071730268315   0.9016265929280587   0.35292301225057904
0.8943733710974386   0.25976047238839683   0.09942746109658186   0.4774609214758912   0.07310813801909873   0.7000022302481936   0.7796642708130705   0.47617723521080674   0.6027819723624176   0.13856418873356813   0.1525850927936481   0.32408810238335034   0.05234507022681615   0.2536669390055239   0.7357845147012521   0.19373174126178613   0.20974064002358683   0.7556066413449952   0.32390704502678314   0.14365518582542655   0.20542094426675217   0.435155924042312   0.4222804520987244   0.7907321735748475   0.31104757316931353   0.17539545165391518   0.32285299100214254   0.31327125209895623   0.2379394351502148   0.4753932214057216   0.543188720189072   0.8370940168881496   0.6351574627877972   0.33682903267215347   0.3906036273954239   0.5130059145047992   0.582812392560981   0.08316209366662959   0.6548191126941719   0.319274173243013   0.37307175253739416   0.3275554523216344   0.3309120676673888   0.17561898741758647   0.167650808270642   0.8923995282793223   0.9086316155686643   0.384886813842739   0.8566032351013285   0.7170040766254072   0.5857786245665219   0.07161556174378272   0.6186637999511136   0.2416108552196856   0.042589904377449826   0.23452154485563323   0.9835063371633165   0.9047818225475321   0.6519862769820259   0.7215156303508341   0.4006939446023355   0.8216197288809025   0.997167164287854   0.4022414571078211
0.027622192064941323   0.49406427655926816   0.6662550966204652   0.22662246969023464   0.8599713837942993   0.6016647482799458   0.7576234810518009   0.8417356558474957   0.00336814869297084   0.8846606716545387   0.17184485648527897   0.770120094103713   0.38470434874185716   0.643049816434853   0.12925495210782917   0.5355985492480797   0.4011980115785406   0.7382679938873209   0.4772686751258033   0.8140829188972456   0.0005040669762051285   0.9166482650064184   0.4801015108379493   0.41184146178942455   0.9728818749112638   0.4225839884471502   0.813846414217484   0.1852189920991899   0.11291049111696448   0.8209192401672044   0.05622293316568322   0.34348333625169425   0.10954234242399363   0.9362585685126659   0.8843780766804042   0.5733632421479813   0.7248379936821365   0.2932087520778128   0.755123124572575   0.03776469289990164   0.32363998210359585   0.5549407581904918   0.2778544494467718   0.22368177400265601   0.3231359151273907   0.6382924931840736   0.7977529386088226   0.8118403122132315   0.35025404021612694   0.21570850473692327   0.9839065243913385   0.6266213201140416   0.23734354909916244   0.3947892645697188   0.9276835912256552   0.28313798386234734   0.1278012066751688   0.458530696057053   0.04330551454525103   0.7097747417143659   0.40296321299303234   0.1653219439792402   0.288182389972676   0.6720100488144644
0.07932323088943646   0.6103811857887483   0.010327940525904147   0.4483282748118083   0.7561873157620457   0.9720886926046748   0.21257500191708162   0.6364879625985769   0.4059332755459188   0.7563801878677515   0.22866847752574312   0.009866642484535233   0.16858972644675635   0.3615909232980327   0.30098488630008785   0.7267286586221879   0.04078851977158755   0.9030602272409798   0.25767937175483685   0.016953916907821925   0.6378253067785552   0.7377382832617395   0.9694969817821608   0.3449438680933576   0.5585020758891188   0.12735709747299123   0.9591690412562567   0.8966155932815493   0.802314760127073   0.15526840486831642   0.7465940393391751   0.26012763068297245   0.39638148458115424   0.39888821700056487   0.517925561813432   0.25026098819843723   0.2277917581343979   0.0372972937025321   0.21694067551334414   0.5235323295762493   0.18700323836281033   0.13423706646155234   0.9592613037585073   0.5065784126684274   0.5491779315842551   0.3964987831998128   0.9897643219763465   0.1616345445750698   0.9906758556951363   0.26914168572682157   0.030595280720089723   0.26501895129352054   0.18836109556806327   0.11387328085850515   0.2840012413809146   0.004891320610548076   0.791979610986909   0.7149850638579403   0.7660756795674826   0.7546303324121109   0.5641878528525112   0.6776877701554082   0.5491350040541385   0.23109800283586154
0.3771846144897008   0.5434507036938558   0.5898737002956311   0.7245195901674342   0.8280066829054458   0.14695192049404307   0.6001093783192847   0.5628850455923644   0.8373308272103094   0.8778102347672215   0.569514097599195   0.2978660942988438   0.6489697316422461   0.7639369539087164   0.2855128562182804   0.2929747736882958   0.8569901206553371   0.04895189005077606   0.5194371766507978   0.5383444412761849   0.2928022678028259   0.37126411989536784   0.9703021725966593   0.30724643844032334   0.9156176533131252   0.8278134162015119   0.3804284723010281   0.5827268482728892   0.08761097040767941   0.6808614957074689   0.7803190939817434   0.01984180268052483   0.25028014319737   0.8030512609402474   0.2108049963825484   0.721975708381681   0.6013104115551239   0.039114307031531036   0.925292140164268   0.42900093469338524   0.7443202908997868   0.990162416980755   0.4058549635134702   0.8906564934172003   0.4515180230969609   0.6188982970853871   0.43555279091681093   0.583410054976877   0.5359003697838357   0.7910848808838752   0.055124318615782805   0.0006832067039877893   0.4482893993761563   0.11022338517640622   0.2748052246340394   0.980841404023463   0.1980092561787863   0.3071721242361588   0.064000228251491   0.25886569564178197   0.5966988446236624   0.2680578172046278   0.138708088087223   0.8298647609483967
0.8523785537238756   0.27789540022387277   0.7328531245737527   0.9392082675311964   0.4008605306269147   0.6589971031384857   0.29730033365694186   0.3557982125543194   0.8649601608430789   0.8679122222546105   0.24217601504115904   0.3551150058503316   0.4166707614669226   0.7576888370782043   0.9673707904071196   0.37427360182686864   0.2186615052881363   0.45051671284204553   0.9033705621556286   0.1154079061850867   0.6219626606644739   0.18245889563741774   0.7646624740684056   0.28554314523668994   0.7695841069405983   0.904563495413545   0.031809349494652854   0.3463348777054936   0.36872357631368363   0.2455663922750593   0.734509015837711   0.9905366651511741   0.5037634154706048   0.37765417002044877   0.49233300079655196   0.6354216593008425   0.0870926540036821   0.6199653329422444   0.5249622103894322   0.2611480574739739   0.8684311487155458   0.1694486201001989   0.6215916482338036   0.14574015128888718   0.24646848805107188   0.9869897244627811   0.856929174165398   0.8601970060521972   0.47688438111047354   0.0824262290492362   0.8251198246707452   0.5138621283467036   0.1081608047967899   0.8368598367741769   0.09061080883303417   0.5233254631955294   0.6043973893261851   0.45920566675372815   0.5982778080364822   0.8879038038946869   0.5173047353225031   0.8392403338114837   0.07331559764704991   0.6267557464207131
0.6488735866069573   0.6697917137112848   0.45172394941324623   0.48101559513182585   0.40240509855588535   0.6828019892485037   0.5947947752478482   0.6208185890796286   0.9255207174454119   0.6003757601992674   0.769674950577103   0.10695646073292502   0.817359912648622   0.7635159234250906   0.6790641417440689   0.5836309975373956   0.21296252332243676   0.3043102566713624   0.08078633370758667   0.6957271936427086   0.6956577879999337   0.4650699228598787   0.00747073606053675   0.06897144722199558   0.046784201392976406   0.7952782091485939   0.5557467866472905   0.5879558520901698   0.644379102837091   0.11247621990009025   0.9609520113994423   0.967137263010541   0.7188583853916792   0.5121004597008229   0.19127706082233922   0.8601808022776161   0.9014984727430573   0.7485845362757323   0.5122129190782704   0.2765498047402205   0.6885359494206205   0.4442742796043699   0.4314265853706837   0.5808226110975119   0.9928781614206869   0.9792043567444911   0.4239558493101469   0.5118511638755163   0.9460939600277104   0.1839261475958973   0.8682090626628565   0.9238953117853466   0.3017148571906194   0.07144992769580702   0.9072570512634142   0.9567580487748055   0.5828564717989402   0.5593494679949842   0.715979990441075   0.09657724649718948   0.6813579990558829   0.8107649317192519   0.2037670713628046   0.820027441756969
0.9928220496352624   0.3664906521148821   0.7723404859921209   0.2392048306594571   0.9999438882145756   0.3872862953703909   0.348384636681974   0.7273536667839408   0.05384992818686518   0.2033601477744936   0.4801755740191176   0.8034583549985942   0.7521350709962458   0.13191022007868658   0.5729185227557034   0.8467003062237887   0.1692785991973056   0.5725607520837024   0.8569385323146285   0.7501230597265992   0.4879206001414227   0.7617958203644505   0.6531714609518239   0.9300956179696303   0.49509855050616025   0.39530516824956835   0.880830974959703   0.6908907873101732   0.4951546622915846   0.008018872879177495   0.5324463382777289   0.9635371205262323   0.44130473410471943   0.804658725104684   0.05227076425861135   0.16007876552763814   0.6891696631084737   0.6727485050259974   0.4793522415029079   0.31337845930384944   0.519891063911168   0.10018775294229496   0.6224137091882794   0.5632553995772502   0.03197046376974541   0.3383919325778445   0.9692422482364554   0.63315978160762   0.5368719132635852   0.9430867643282761   0.08841127327675252   0.9422689942974469   0.04171725097200054   0.9350678914490986   0.5559649349990236   0.9787318737712146   0.600412516867281   0.13040916634441477   0.5036941707404122   0.8186531082435765   0.9112428537588074   0.4576606613184174   0.02434192923750432   0.505274648939727
0.39135178984763935   0.3574729083761225   0.4019282200492249   0.9420192493624767   0.3593813260778939   0.01908097579827796   0.43268597181276947   0.30885946775485673   0.8225094128143088   0.07599421147000182   0.34427469853601694   0.3665904734574098   0.7807921618423083   0.14092632002090316   0.7883097635369933   0.38785859968619524   0.18037964497502715   0.01051715367648841   0.2846155927965811   0.5692054914426188   0.2691367912162197   0.552856492358071   0.2602736635590768   0.06393084250289174   0.8777850013685804   0.1953835839819485   0.8583454435098519   0.12191159314041498   0.5184036752906864   0.17630260818367052   0.42565947169708246   0.8130521253855583   0.6958942624763776   0.10030839671366872   0.08138477316106552   0.44646165192814846   0.9151021006340695   0.9593820766927655   0.2930750096240722   0.058603052241953266   0.7347224556590424   0.9488649230162771   0.008459416827491056   0.4893975607993345   0.4655856644428226   0.3960084306582062   0.7481857532684143   0.4254667182964428   0.5878006630742422   0.20062484667625766   0.8898403097585624   0.3035551251560278   0.06939698778355578   0.024322238492587134   0.46418083806148   0.4905029997704695   0.3735027253071781   0.9240138417789184   0.3827960649004144   0.04404134784232103   0.45840062467310866   0.9646317650861529   0.08972105527634225   0.9854382956003678
0.7236781690140663   0.015766842069875723   0.08126163844885119   0.4960407348010332   0.2580925045712437   0.6197584114116695   0.33307588518043696   0.07057401650459048   0.6702918414970015   0.4191335647354119   0.4432355754218746   0.7670188913485627   0.6008948537134458   0.3948113262428248   0.9790547373603946   0.2765158915780932   0.22739212840626763   0.47079748446390635   0.5962586724599802   0.23247454373577217   0.7689915037331589   0.5061657193777535   0.506537617183638   0.2470362481354044   0.04531333471909268   0.49039887730787773   0.42527597873478673   0.7509955133343712   0.7872208301478489   0.8706404658962081   0.0922000935543498   0.6804214968297807   0.11692898865084747   0.4515069011607963   0.6489645181324752   0.913402605481218   0.5160341349374018   0.056695574917971545   0.6699097807720806   0.6368867139031248   0.28864200653113414   0.5858980904540652   0.07365110831210045   0.4044121701673526   0.5196505027979751   0.07973237107631173   0.5671134911284625   0.1573759220319482   0.47433716807888243   0.589333493768434   0.14183751239367579   0.406380408697577   0.6871163379310335   0.7186930278722258   0.049637418839325965   0.7259589118677964   0.570187349280186   0.2671861267114295   0.40067290070685074   0.8125563063865784   0.05415321434278428   0.21049055179345794   0.7307631199347701   0.17566959248345362
0.7655112078116502   0.6245924613393927   0.6571120116226696   0.7712574223161011   0.24586070501367502   0.544860090263081   0.0899985204942071   0.6138815002841528   0.7715235369347926   0.955526596494647   0.9481610081005314   0.20750109158657576   0.08440719900375906   0.23683356862242122   0.8985235892612053   0.4815421797187794   0.514219849723573   0.9696474419109917   0.49785068855435466   0.668985873332201   0.46006663538078874   0.7591568901175338   0.7670875686195846   0.4933162808487474   0.6945554275691386   0.1345644287781411   0.10997555699691496   0.7220588585326464   0.4486947225554636   0.5897043385150601   0.019977036502707844   0.1081773582484936   0.677171185620671   0.6341777420204131   0.0718160284021765   0.9006762666619178   0.592763986616912   0.39734417339799183   0.17329243914097114   0.4191340869431384   0.0785441368933389   0.4276967314870001   0.6754417505866165   0.7501482136109374   0.6184775015125501   0.6685398413694663   0.9083541819670319   0.25683193276218996   0.9239220739434115   0.5339754125913252   0.7983786249701169   0.5347730742295436   0.47522735138794797   0.9442710740762651   0.7784015884674091   0.42659571598104995   0.7980561657672769   0.31009333205585204   0.7065855600652327   0.5259194493191321   0.205292179150365   0.9127491586578602   0.5332931209242615   0.10678536237599373
0.12674804225702607   0.4850524271708601   0.857851370337645   0.35663714876505637   0.508270540744476   0.8165125858013939   0.949497188370613   0.09980521600286636   0.5843484668010643   0.2825371732100686   0.15111856340049612   0.5650321417733228   0.10912111541311643   0.3382660991338035   0.37271697493308703   0.13843642579227283   0.31106494964583953   0.028172767077951473   0.6661314148678544   0.6125169764731406   0.10577277049547454   0.11542360842009126   0.13283829394359295   0.505731614097147   0.9790247282384484   0.6303711812492312   0.27498692360594795   0.14909446533209061   0.4707541874939725   0.8138585954478373   0.32548973523533486   0.049289249329224245   0.8864057206929081   0.5313214222377687   0.17437117183483877   0.48425710755590146   0.7772846052797917   0.1930553231039652   0.8016541969017518   0.3458206817636286   0.4662196556339522   0.1648825560260137   0.13552278203389737   0.7333037052904879   0.36044688513847767   0.04945894760592245   0.0026844880903044146   0.22757209119334101   0.3814221569000292   0.41908776635669126   0.7276975644843564   0.07847762586125041   0.9106679694060567   0.605229170908854   0.40220782924902154   0.029188376532026168   0.02426224871314852   0.07390774867108525   0.2278366574141828   0.5449312689761248   0.24697764343335682   0.8808524255671201   0.426182460512431   0.19911058721249608
0.7807579877994046   0.7159698695411063   0.2906596784785337   0.46580688192200814   0.42031110266092697   0.6665109219351839   0.2879751903882293   0.23823479072866713   0.03888894576089777   0.24742315557849262   0.5602776259038729   0.1597571648674167   0.12822097635484112   0.6421939846696386   0.15806979665485124   0.13056878833539054   0.10395872764169259   0.5682862359985534   0.9302331392406684   0.5856375193592658   0.8569810842083357   0.6874338104314334   0.5040506787282374   0.38652693214676975   0.07622309640893114   0.9714639408903271   0.21339100024970373   0.9207200502247616   0.6559119937480041   0.3049530189551431   0.9254158098614744   0.6824852594960945   0.6170230479871064   0.0575298633766505   0.3651381839576016   0.5227280946286778   0.4888020716322653   0.41533587870701183   0.20706838730275037   0.3921593062932872   0.38484334399057274   0.8470496427084584   0.27683524806208193   0.8065217869340214   0.527862259782237   0.15961583227702508   0.7727845693338445   0.4199948547872517   0.45163916337330584   0.18815189138669808   0.5593935690841408   0.49927480456249007   0.7957271696253017   0.8831988724315549   0.6339777592226663   0.8167895450663956   0.17870412163819524   0.8256690090549045   0.26883957526506475   0.2940614504377178   0.68990205000593   0.41033313034789265   0.06177118796231434   0.9019021441444306
0.30505870601535723   0.5632834876394341   0.7849359399002324   0.09538035721040913   0.7771964462331202   0.4036676553624091   0.012151370566387869   0.6753855024231574   0.32555728285981445   0.215515763975711   0.45275780148224704   0.17611069786066738   0.5298301132345128   0.33231689154415606   0.8187800422595807   0.3593211527942718   0.3511259915963176   0.5066478824892515   0.5499404669945159   0.06525970235655403   0.6612239415903877   0.09631475214135893   0.48816927903220164   0.16335755821212347   0.3561652355750304   0.5330312645019247   0.7032333391319693   0.06797720100171434   0.5789687893419101   0.12936360913951564   0.6910819685655814   0.39259169857855686   0.2534115064820957   0.9138478451638047   0.23832416708333432   0.2164810007178895   0.7235813932475829   0.5815309536196486   0.4195441248237536   0.8571598479236177   0.37245540165126534   0.07488307113039705   0.8696036578292377   0.7919001455670637   0.7112314600608777   0.9785683189890381   0.381434378797036   0.6285425873549402   0.3550662244858473   0.4455370544871134   0.6782010396650667   0.5605653863532258   0.7760974351439371   0.3161734453475977   0.9871190710994854   0.16797368777466892   0.5226859286618415   0.4023256001837931   0.7487949040161511   0.9514926870567795   0.7991045354142586   0.8207946465641445   0.3292507791923975   0.09433283913316177
0.42664913376299324   0.7459115754337474   0.4596471213631598   0.30243269356609814   0.7154176737021156   0.7673432564447092   0.07821274256612384   0.673890106211158   0.36035144921626827   0.3218062019575959   0.4000117029010571   0.11332471985793215   0.5842540140723311   0.005632756609998214   0.4128926318015717   0.9453510320832632   0.061568085410489644   0.6033071564262051   0.6640977277854206   0.9938583450264837   0.26246354999623106   0.7825125098620607   0.3348469485930232   0.899525505893322   0.8358144162332378   0.03660093442831327   0.8751998272298633   0.5970928123272239   0.12039674253112223   0.26925767798360395   0.7969870846637396   0.9232027061160659   0.7600452933148539   0.9474514760260081   0.39697538176268243   0.8098779862581338   0.17579127924252283   0.9418187194160098   0.9840827499611107   0.8645269541748706   0.11422319383203319   0.33851156298980467   0.3199850221756901   0.8706686091483867   0.8517596438358022   0.555999053127744   0.9851380735826669   0.9711431032550648   0.015945227602564345   0.5193981186994308   0.1099382463528035   0.3740502909278409   0.8955484850714421   0.25014044071582675   0.312951161689064   0.450847584811775   0.13550319175658818   0.3026889646898187   0.9159757799263816   0.6409695985536412   0.9597119125140653   0.3608702452738089   0.9318930299652708   0.7764426443787708
0.8454887186820321   0.022358682284004196   0.6119080077895808   0.9057740352303839   0.99372907484623   0.46635962915626017   0.626769934206914   0.9346309319753191   0.9777838472436656   0.9469615104568294   0.5168316878541104   0.5605806410474782   0.08223536217222352   0.6968210697410027   0.20388052616504643   0.1097330562357032   0.9467321704156354   0.394132105051184   0.2879047462386649   0.46876345768206196   0.98702025790157   0.033261859777375107   0.35601171627339406   0.6923208133032912   0.1415315392195379   0.01090317749337091   0.7441037084838132   0.7865467780729073   0.1478024643733079   0.5445435483371107   0.11733377427689934   0.8519158460975882   0.17001861712964225   0.5975820378802813   0.6005020864227889   0.2913352050501099   0.08778325495741873   0.9007609681392785   0.3966215602577425   0.1816021488144067   0.14105108454178336   0.5066288630880945   0.1087168140190776   0.7128386911323448   0.15403082664021334   0.47336700331071946   0.7527050977456836   0.02051787782905354   0.012499287420675444   0.4624638258173485   0.008601389261870306   0.23397109975614624   0.8646968230473675   0.9179202774802379   0.891267614984971   0.38205525365855814   0.6946782059177253   0.32033823959995655   0.2907655285621821   0.0907200486084482   0.6068949509603065   0.419577271460678   0.8941439683044395   0.9091178997940415
0.4658438664185232   0.9129484083725835   0.7854271542853619   0.19627920866169674   0.3118130397783099   0.439581405061864   0.032722056539678405   0.1757613308326432   0.2993137523576344   0.9771175792445155   0.024120667277808098   0.941790231076497   0.43461692931026685   0.05919730176427766   0.13285305229283711   0.5597349774179389   0.7399387233925415   0.7388590621643211   0.8420875237306551   0.4690149288094906   0.133043772432235   0.3192817907036431   0.9479435554262156   0.5598970290154491   0.6671999060137118   0.4063333823310596   0.16251640114085356   0.36361782035375234   0.355386866235402   0.9667519772691956   0.12979434460117514   0.18785648952110917   0.05607311387776757   0.9896343980246801   0.10567367732336705   0.24606625844461222   0.6214561845675007   0.9304370962604025   0.9728206250305299   0.6863312810266734   0.8815174611749591   0.19157803409608135   0.13073310129987484   0.21731635221718282   0.7484736887427241   0.8722962433924383   0.18278954587365934   0.6574193232017337   0.0812737827290123   0.4659628610613787   0.020273144732805778   0.29380150284798134   0.7258869164936104   0.4992108837921831   0.8904788001316306   0.10594501332687216   0.6698138026158428   0.5095764857675029   0.7848051228082635   0.85987875488226   0.04835761804834205   0.5791393895071005   0.8119844977777336   0.17354747385558653
0.1668401568733829   0.38756135541101916   0.6812513964778588   0.9562311216384037   0.4183664681306588   0.5152651120185809   0.4984618506041995   0.29881179843667   0.3370926854016465   0.04930225095720225   0.4781887058713937   0.005010295588688679   0.6112057689080362   0.5500913671650192   0.5877099057397631   0.8990652822618165   0.9413919662921935   0.0405148813975162   0.8029047829314995   0.03918652737955658   0.8930343482438514   0.46137549189041566   0.9909202851537658   0.8656390535239701   0.7261941913704685   0.0738141364793965   0.30966888867590703   0.9094079318855663   0.30782772323980967   0.5585490244608156   0.8112070380717075   0.6105961334488963   0.9707350378381632   0.5092467735036134   0.3330183322003138   0.6055858378602077   0.35952926893012693   0.9591554063385942   0.7453084264605506   0.7065205555983911   0.4181373026379335   0.918640524941078   0.9424036435290511   0.6673340282188346   0.525102954394082   0.4572650330506623   0.9514833583752853   0.8016949746948645   0.7989087630236137   0.3834508965712658   0.6418144696993783   0.8922870428092982   0.49108103978380396   0.8249018721104502   0.8306074316276708   0.2816909093604018   0.5203460019456408   0.3156550986068369   0.497589099427357   0.6761050715001942   0.16081673301551389   0.35649969226824274   0.7522806729668063   0.9695845159018031
0.7426794303775804   0.43785916732716473   0.8098770294377552   0.30225048768296847   0.21757647598349827   0.9805941342765024   0.8583936710624699   0.500555512988104   0.41866771295988464   0.5971432377052367   0.21657920136309158   0.6082684701788058   0.9275866731760807   0.7722413655947864   0.3859717697354208   0.326577560818404   0.40724067123043983   0.4565862669879496   0.8883826703080637   0.6504724893182099   0.24642393821492595   0.10008657471970683   0.13610199734125736   0.6808879734164068   0.5037445078373456   0.662227407392542   0.32622496790350214   0.37863748573343836   0.28616803185384726   0.6816332731160396   0.46783129684103225   0.8780819727453344   0.8675003188939626   0.08449003541080298   0.25125209547794064   0.2698135025665286   0.9399136457178819   0.3122486698160165   0.8652803257425199   0.9432359417481246   0.5326729744874421   0.8556624028280669   0.9768976554344562   0.29276345242991475   0.2862490362725162   0.7555758281083601   0.8407956580931988   0.6118754790135079   0.7825045284351706   0.09334842071581806   0.5145706901896966   0.23323799328006956   0.49633649658132334   0.41171514759977845   0.046739393348664386   0.35515602053473516   0.6288361776873608   0.32722511218897543   0.7954872978707237   0.08534251796820655   0.6889225319694787   0.014976442372958913   0.9302069721282038   0.14210657622008196
0.15624955748203664   0.15931403954489193   0.9533093166937477   0.8493431237901672   0.8700005212095204   0.40373821143653177   0.11251365860054893   0.2374676447766593   0.08749599277434984   0.3103897907207137   0.5979429684108523   0.0042296514965897355   0.5911594961930264   0.8986746431209353   0.5512035750621879   0.6490736309618546   0.9623233185056658   0.5714495309319598   0.7557162771914642   0.5637311129936481   0.273400786536187   0.5564730885590009   0.8255093050632604   0.4216245367735661   0.11715122905415033   0.39715904901410903   0.8721999883695126   0.5722814129833989   0.24715070784462986   0.9934208375775773   0.7596863297689637   0.3348137682067396   0.15965471507028   0.6830310468568634   0.16174336135811138   0.33058411671014987   0.5684952188772535   0.7843564037359282   0.6105397862959234   0.6815104857482952   0.6061719003715877   0.21290687280396833   0.8548235091044593   0.11777937275464721   0.3327711138354008   0.6564337842449673   0.02931420404119893   0.6961548359810812   0.21561988478125046   0.25927473523085837   0.15711421567168632   0.12387342299768227   0.9684691769366206   0.26585389765328116   0.3974278859027226   0.7890596547909426   0.8088144618663405   0.5828228507964177   0.23568452454461125   0.45847553808079283   0.24031924298908705   0.7984664470604895   0.6251447382486878   0.7769650523324976
0.6341473426174993   0.5855595742565212   0.7703212291442285   0.6591856795778503   0.30137622878209847   0.9291257900115537   0.7410070251030296   0.9630308435967693   0.08575634400084801   0.6698510547806954   0.5838928094313433   0.8391574205990869   0.1172871670642274   0.4039971571274142   0.18646492352862065   0.05009776580814428   0.30847270519788683   0.8211743063309965   0.9507803989840095   0.5916222277273514   0.06815346220879974   0.022707859270507065   0.32563566073532163   0.8146571753948538   0.4340061195913005   0.43714828501398595   0.5553144315910931   0.1554714958170035   0.13262989080920198   0.5080224950024321   0.8143074064880635   0.1924406522202343   0.04687354680835396   0.8381714402217368   0.23041459705672027   0.35328323162114733   0.9295863797441266   0.4341742830943226   0.04394967352809961   0.30318546581300304   0.6211136745462398   0.6129999767633261   0.0931692745440902   0.7115632380856516   0.55296021233744   0.590292117492819   0.7675336138087686   0.8969060626907978   0.11895409274613955   0.15314383247883306   0.21221918221767547   0.7414345668737942   0.9863242019369376   0.6451213374764009   0.39791177572961195   0.54899391465356   0.9394506551285836   0.806949897254664   0.16749717867289168   0.19571068303241257   0.009864275384457047   0.3727756141603415   0.12354750514479207   0.8925252172194096
0.3887506008382173   0.7597756373970154   0.03037823060070187   0.18096197913375794   0.8357903885007772   0.1694835199041964   0.2628446167919333   0.2840559164429602   0.7168362957546377   0.016339687425363323   0.05062543457425785   0.542621349569166   0.7305120938177001   0.3712183499489624   0.6527136588446459   0.9936274349156061   0.7910614386891165   0.5642684526942984   0.4852164801717542   0.7979167518831936   0.7811971633046595   0.19149283853395688   0.36166897502696216   0.905391534663784   0.3924465624664422   0.43171720113694145   0.33129074442626033   0.7244295555300261   0.5566561739656649   0.26223368123274504   0.06844612763432702   0.44037363908706584   0.8398198782110272   0.24589399380738175   0.017820693060069167   0.8977522895178999   0.10930778439332706   0.8746756438584193   0.36510703421542323   0.9041248546022937   0.3182463457042105   0.31040719116412097   0.879890554043669   0.10620810271910022   0.537049182399551   0.11891435263016412   0.5182215790167068   0.20081656805531625   0.14460261993310886   0.6871971514932227   0.18693083459044652   0.4763870125252902   0.5879464459674439   0.4249634702604776   0.1184847069561195   0.03601337343822436   0.7481265677564167   0.17906947645309582   0.10066401389605033   0.13826108392032452   0.6388187833630896   0.3043938325946765   0.735556979680627   0.2341362293180308
0.3205724376588791   0.9939866414305555   0.855666425636958   0.12792812659893057   0.7835232552593281   0.8750722888003915   0.33744484662025126   0.9271115585436143   0.6389206353262192   0.18787513730716876   0.15051401202980474   0.4507245460183241   0.0509741893587753   0.7629116670466912   0.03202930507368527   0.41471117258009976   0.30284762160235856   0.5838421905935953   0.9313652911776349   0.2764500886597752   0.664028838239269   0.2794483579989189   0.19580831149700786   0.042313859341744434   0.3434564005803898   0.28546171656836333   0.3401418858600498   0.9143857327428139   0.5599331453210616   0.41038942776797194   0.0026970392397985227   0.9872741741991996   0.9210125099948424   0.22251429046080315   0.8521830272099937   0.5365496281808755   0.8700383206360671   0.45960262341411195   0.8201537221363085   0.12183845560077568   0.5671906990337086   0.8757604328205166   0.8887884309586735   0.8453883669410005   0.9031618607944397   0.5963120748215978   0.6929801194616657   0.803074507599256   0.5597054602140499   0.3108503582532344   0.3528382336016159   0.8886887748564422   0.9997723148929882   0.9004609304852624   0.3501411943618174   0.9014146006572427   0.07875980489814578   0.6779466400244594   0.4979581671518236   0.3648649724763672   0.20872148426207862   0.21834401661034736   0.6778044450155152   0.2430265168755915
0.64153078522837   0.3425835837898307   0.7890160140568415   0.397638149934591   0.7383689244339303   0.746271508968233   0.09603589459517586   0.594563642335335   0.1786634642198804   0.4354211507149986   0.74319766099356   0.7058748674788928   0.17889114932689218   0.5349602202297361   0.39305646663174254   0.8044602668216502   0.10013134442874638   0.8570135802052767   0.8950982994799189   0.43959529434528305   0.8914098601666678   0.6386695635949294   0.2172938544644038   0.19656877746969156   0.24987907493829772   0.2960859798050987   0.4282778404075622   0.7989306275351005   0.5115101505043674   0.5498144708368657   0.33224194581238636   0.2043669851997655   0.332846686284487   0.11439332012186709   0.5890442848188264   0.4984921177208727   0.1539555369575948   0.579433099892131   0.19598781818708386   0.6940318508992225   0.05382419252884842   0.7224195196868543   0.30088951870716496   0.25443655655393943   0.16241433236218067   0.08374995609192476   0.08359566424276116   0.05786777908424785   0.912535257423883   0.787663976286826   0.6553178238351989   0.2589371515491473   0.40102510691951554   0.23784950544996036   0.32307587802281257   0.05457016634938181   0.06817842063502855   0.12345618532809328   0.7340315932039861   0.5560780486285092   0.9142228836774338   0.5440230854359623   0.5380437750169023   0.8620461977292867
0.8603986911485854   0.8216035657491081   0.23715425630973733   0.6076096411753472   0.6979843587864046   0.7378536096571834   0.15355859206697617   0.5497418620910994   0.7854491013625217   0.9501896333703572   0.49824076823177726   0.29080471054195206   0.3844239944430062   0.7123401279203969   0.17516489020896467   0.23623454419257028   0.31624557380797763   0.5888839425923036   0.4411332970049785   0.6801564955640611   0.4020226901305439   0.044860857156341326   0.9030895219880762   0.8181102978347745   0.5416239989819586   0.22325729140723322   0.6659352656783389   0.21050065665942722   0.8436396401955539   0.4854036817500499   0.5123766736113627   0.6607587945683278   0.05819053883303224   0.5352140483796926   0.014135905379585511   0.3699540840263757   0.673766544390026   0.8228739204592957   0.8389710151706209   0.13371953983380544   0.3575209705820484   0.23398997786699208   0.39783771816564234   0.45356304426974425   0.9554982804515045   0.18912912071065074   0.49474819617756605   0.6354527464349699   0.4138742814695459   0.9658718293034175   0.8288129304992271   0.4249520897755426   0.5702346412739919   0.48046814755336764   0.3164362568878644   0.7641932952072148   0.5120441024409597   0.9452540991736751   0.3023003515082789   0.3942392111808391   0.8382775580509336   0.12238017871437934   0.46332933633765805   0.2605196713470337
0.4807565874688852   0.8883902008473873   0.06549161817201574   0.8069566270772894   0.5252583070173807   0.6992610801367365   0.5707434219944497   0.17150388064231958   0.11138402554783483   0.733389250833319   0.7419304914952225   0.746551790866777   0.5411493842738428   0.2529211032799513   0.42549423460735813   0.9823584956595622   0.029105281832883183   0.3076670041062763   0.12319388309907923   0.5881192844787231   0.19082772378194954   0.18528682539189692   0.6598645467614211   0.3275996131316894   0.7100711363130643   0.29689662454450966   0.5943729285894055   0.5206429860544001   0.18481282929568355   0.5976355444077732   0.0236295065949558   0.34913910541208043   0.07342880374784871   0.8642462935744543   0.2816990150997333   0.6025873145453035   0.5322794194740058   0.6113251902945029   0.8562047804923751   0.6202288188857412   0.5031741376411226   0.30365818618822665   0.733010897393296   0.032109534407018164   0.3123464138591731   0.11837136079632969   0.07314635063187473   0.7045099212753287   0.6022752775461089   0.82147473625182   0.47877342204246925   0.1838669352209287   0.4174624482504253   0.22383919184404683   0.4551439154475135   0.8347278298088483   0.34403364450257656   0.3595928982695926   0.17344490034778018   0.23214051526354482   0.8117542250285708   0.7482677079750897   0.317240119855405   0.6119116963778036
0.3085800873874481   0.4446095217868631   0.5842292224621091   0.5798021619707854   0.996233673528275   0.3262381609905334   0.5110828718302344   0.8752922406954566   0.39395839598216614   0.5047634247387134   0.0323094497877651   0.691425305474528   0.9764959477317409   0.28092423289466656   0.5771655343402516   0.8566974756656797   0.6324623032291643   0.9213313346250739   0.4037206339924715   0.6245569604021348   0.8207080782005935   0.1730636266499842   0.08648051413706646   0.012645264024331275   0.5121279908131454   0.7284541048631211   0.5022512916749574   0.43284310205354587   0.5158943172848705   0.4022159438725877   0.991168419844723   0.5575508613580892   0.12193592130270432   0.8974525191338744   0.9588589700569579   0.8661255558835612   0.14543997357096344   0.6165282862392077   0.3816934357167063   0.009428080217881569   0.5129776703417991   0.6951969516141339   0.9779728017242348   0.38487111981574673   0.6922695921412055   0.5221333249641497   0.8914922875871684   0.3722258557914154   0.18014160132806006   0.7936792201010285   0.38924099591221095   0.9393827537378696   0.6642472840431896   0.39146327622844085   0.39807257606748797   0.3818318923797804   0.5423113627404853   0.49401075709456654   0.43921360601053006   0.5157063364962191   0.3968713891695218   0.8774824708553588   0.057520170293823766   0.5062782562783376
0.8838937188277227   0.18228551924122494   0.07954736856958897   0.12140713646259084   0.19162412668651718   0.6601521942770753   0.18805508098242063   0.7491812806711754   0.0114825253584571   0.8664729741760467   0.7988140850702097   0.8097985269333058   0.3472352413152675   0.4750096979476059   0.4007415090027217   0.42796663455352546   0.8049238785747822   0.9809989408530394   0.9615279029921917   0.9122602980573064   0.4080524894052604   0.1035164699976806   0.904007732698368   0.40598204177896874   0.5241587705775377   0.9212309507564557   0.824460364128779   0.2845749053163779   0.33253464389102055   0.2610787564793804   0.6364052831463584   0.5353936246452025   0.32105211853256344   0.39460578230333365   0.8375911980761487   0.7255950977118967   0.9738168772172959   0.9195960843557277   0.4368496890734269   0.2976284631583712   0.16889299864251367   0.9385971435026883   0.4753217860812352   0.3853681651010649   0.7608405092372532   0.8350806735050077   0.5713140533828673   0.9793861233220962   0.23668173865971556   0.913849722748552   0.7468536892540883   0.6948112180057183   0.904147094768695   0.6527709662691717   0.11044840610773   0.15941759336051584   0.5830949762361316   0.25816518396583804   0.27285720803158137   0.43382249564861913   0.6092780990188357   0.33856909961011034   0.8360075189581544   0.13619403249024792
0.440385100376322   0.399971956107422   0.36068573287691924   0.750825867389183   0.6795445911390687   0.5648912826024143   0.789371679494052   0.7714397440670868   0.4428628524793532   0.6510415598538621   0.04251799023996359   0.07662852606136847   0.5387157577106582   0.9982705935846905   0.9320695841322336   0.9172109327008526   0.9556207814745266   0.7401054096188524   0.6592123761006522   0.4833884370522335   0.3463426824556909   0.40153631000874207   0.8232048571424978   0.3471944045619856   0.9059575820793688   0.0015643539013200775   0.46251912426557856   0.5963685371728026   0.2264129909403001   0.4366730712989058   0.6731474447715267   0.8249287931057159   0.7835501384609469   0.7856315114450436   0.630629454531563   0.7483002670443474   0.24483438075028877   0.7873609178603532   0.6985598703993294   0.8310893343434947   0.2892135992757622   0.04725550824150077   0.03934749429867725   0.34770089729126125   0.9428709168200713   0.6457191982327587   0.21614263715617948   0.0005064927292756467   0.03691333474070247   0.6441548443314387   0.7536235128906009   0.404137955556473   0.8105003438004024   0.2074817730325328   0.08047606811907429   0.5792091624507573   0.026950205339455444   0.4218502615874891   0.44984661358751127   0.8309088954064099   0.7821158245891667   0.634489343727136   0.7512867431881818   0.9998195610629151
0.4929022253134045   0.5872338354856351   0.7119392488895046   0.652118663771654   0.5500313084933331   0.9415146372528764   0.49579661173332507   0.6516121710423782   0.5131179737526307   0.2973597929214378   0.7421730988427241   0.24747421548590523   0.7026176299522283   0.08987801988890506   0.6616970307236498   0.668265053035148   0.6756674246127728   0.6680277583014159   0.21185041713613859   0.8373561576287382   0.8935516000236062   0.03353841457427998   0.46056367394795683   0.837536596565823   0.40064937471020173   0.4463045790886448   0.7486244250584523   0.18541793279416907   0.8506180662168685   0.5047899418357683   0.2528278133251272   0.5338057617517907   0.3375000924642379   0.20743014891433048   0.5106547144824031   0.28633154626588553   0.6348824625120095   0.11755212902542542   0.8489576837587532   0.6180664932307376   0.9592150378992367   0.44952437072400947   0.6371072666226146   0.7807103356019994   0.0656634378756305   0.4159859561497295   0.17654359267465786   0.9431737390361764   0.6650140631654288   0.9696813770610847   0.4279191676162056   0.7577558062420073   0.8143959969485602   0.4648914352253164   0.17509135429107836   0.22395004449021658   0.47689590448432234   0.2574612863109859   0.6644366398086753   0.937618498224331   0.8420134419723128   0.1399091572855605   0.815478956049922   0.3195520049935935
0.8827984040730761   0.690384786561551   0.17837168942730738   0.5388416693915941   0.8171349661974456   0.2743988304118215   0.0018280967526495382   0.5956679303554177   0.1521209030320168   0.30471745335073674   0.573908929136444   0.8379121241134103   0.33772490608345657   0.8398260181254203   0.3988175748453656   0.6139620796231937   0.8608290015991342   0.5823647318144345   0.7343809350366903   0.6763435813988627   0.018815559626821438   0.44245557452887396   0.9189019789867683   0.35679157640526926   0.13601715555374533   0.752070787967323   0.7405302895594609   0.8179499070136752   0.31888218935629975   0.4776719575555015   0.7387021928068114   0.22228197665825755   0.16676128632428291   0.17295450420476471   0.1647932636703674   0.38436985254484723   0.8290363802408264   0.33312848607934437   0.7659756888250018   0.7704077729216535   0.9682073786416922   0.7507637542649099   0.03159475378831148   0.0940641915227908   0.9493918190148707   0.3083081797360359   0.1126927748015432   0.7372726151175215   0.8133746634611253   0.5562373917687129   0.37216248524208234   0.9193227081038464   0.4944924741048256   0.07856543421321145   0.633460292435271   0.6970407314455889   0.32773118778054267   0.9056109300084467   0.46866702876490357   0.3126708789007416   0.49869480753971634   0.5724824439291024   0.7026913399399018   0.5422631059790881
0.5304874288980242   0.8217186896641925   0.6710965861515903   0.4481989144562973   0.5810956098831536   0.5134105099281566   0.5584038113500471   0.7109262993387757   0.7677209464220281   0.9571731181594436   0.1862413261079648   0.7916035912349293   0.2732284723172026   0.8786076839462321   0.5527810336726938   0.0945628597893405   0.9454972845366599   0.9729967539377854   0.08411400490779022   0.7818919808885989   0.44680247699694353   0.4005143100086831   0.3814226649678884   0.23962887490951085   0.9163150480989193   0.5787956203444906   0.7103260788162981   0.7914299604532136   0.3352194382157658   0.06538511041633402   0.151922267466251   0.08050366111443788   0.5674984917937376   0.10821199225689039   0.9656809413582862   0.28890006987950856   0.29427001947653497   0.22960430831065823   0.4128999076855924   0.19433721009016805   0.3487727349398751   0.2566075543728728   0.3287859027778022   0.4124452292015691   0.9019702579429315   0.8560932443641898   0.9473632378099137   0.17281635429205827   0.9856552098440122   0.27729762401969915   0.23703715899361563   0.3813863938388447   0.6504357716282464   0.2119125136033651   0.08511489152736464   0.3008827327244068   0.08293727983450885   0.10370052134647471   0.11943395016907843   0.011982662844898278   0.7886672603579739   0.8740962130358165   0.7065340424834861   0.8176454527547302
0.43989452541809876   0.6174886586629437   0.3777481397056838   0.4052002235531611   0.5379242674751672   0.761395414298754   0.4303849018957701   0.23238386926110283   0.5522690576311551   0.48409779027905486   0.19334774290215445   0.8509974754222581   0.9018332860029086   0.27218527667568976   0.1082328513747898   0.5501147426978513   0.8188960061683997   0.16848475532921503   0.9887989012057113   0.5381320798529531   0.03022874581042591   0.29438854229339856   0.28226485872222534   0.7204866270982228   0.5903342203923271   0.6768998836304548   0.9045167190165415   0.3152864035450617   0.052409952917159885   0.9155044693317008   0.4741318171207714   0.08290253428395886   0.5001408952860048   0.43140667905264596   0.28078407421861695   0.23190505886170074   0.5983076092830962   0.15922140237695623   0.17255122284382718   0.6817903161638494   0.7794116031146965   0.9907366470477412   0.18375232163811578   0.1436582363108964   0.7491828573042705   0.6963481047543426   0.9014874629158904   0.4231716092126736   0.1588486369119434   0.019448221123887798   0.9969707438993489   0.10788520566761191   0.10643868399478351   0.10394375179218696   0.5228389267785775   0.024982671383653048   0.6062977887087787   0.672537072739541   0.2420548525599605   0.7930776125219523   0.007990179425682453   0.5133156703625847   0.06950362971613334   0.1112872963581029
0.22857857631098602   0.5225790233148436   0.8857513080780176   0.9676290600472065   0.47939571900671546   0.8262309185605009   0.9842638451621272   0.5444574508345329   0.32054708209477206   0.8067826974366131   0.9872931012627782   0.436572245166921   0.21410839809998858   0.7028389456444262   0.46445417448420073   0.411589573783268   0.6078106093912099   0.03030187290488521   0.22239932192424022   0.6185119612613157   0.5998204299655274   0.5169862025423004   0.15289569220810686   0.5072246649032127   0.37124185365454143   0.9944071792274569   0.2671443841300893   0.5395956048560062   0.8918461346478259   0.16817626066695593   0.28288053896796217   0.9951381540214733   0.5712990525530539   0.3613935632303428   0.2955874377051839   0.5585659088545523   0.3571906544530653   0.6585546175859166   0.8311332632209832   0.1469763350712843   0.7493800450618554   0.6282527446810314   0.608733941296743   0.5284643738099687   0.14955961509632798   0.11126654213873095   0.4558382490886361   0.021239708906755903   0.7783177614417865   0.11685936291127406   0.18869386495854684   0.4816441040507497   0.8864716267939606   0.9486831022443182   0.9058133259905846   0.4865059500292764   0.3151725742409067   0.5872895390139753   0.6102258882854007   0.9279400411747241   0.9579819197878414   0.9287349214280587   0.7790926250644175   0.7809637061034398
0.208601874725986   0.3004821767470273   0.17035868376767452   0.25249933229347116   0.05904225962965801   0.18921563460829638   0.7145204346790384   0.23125962338671524   0.2807244981878715   0.07235627169702231   0.5258265697204916   0.7496155193359656   0.39425287139391085   0.12367316945270418   0.6200132437299068   0.26310956930668916   0.07908029715300414   0.5363836304387288   0.009787355444506164   0.3351695281319651   0.12109837736516274   0.6076487090106701   0.23069473038008867   0.5542058220285253   0.9124965026391767   0.30716653226364277   0.060336046612414145   0.30170648973505415   0.8534542430095188   0.11795089765534639   0.3458156119333758   0.07044686634833894   0.5727297448216473   0.04559462595832407   0.8199890422128843   0.32083134701237337   0.1784768734277364   0.9219214565056199   0.19997579848297733   0.057721777705684194   0.09939657627473227   0.3855378260668911   0.19018844303847116   0.7225522495737191   0.9782981989095695   0.777889117056221   0.9594937126583825   0.1683464275451938   0.06580169627039278   0.47072258479257817   0.8991576660459684   0.8666399378101396   0.21234745326087404   0.3527716871372318   0.5533420541125926   0.7961930714618007   0.6396177084392267   0.3071770611789077   0.7333530118997084   0.4753617244494273   0.46114083501149034   0.3852556046732878   0.533377213416731   0.4176399467437431
0.3617442587367581   0.9997177786063968   0.3431887703782599   0.695087697170024   0.38344605982718855   0.22182866155017583   0.3836950577198774   0.5267412696248303   0.31764436355679576   0.7511060767575977   0.484537391673909   0.6601013318146906   0.10529691029592173   0.3983343896203659   0.9311953375613164   0.8639082603528899   0.465679201856695   0.09115732844145817   0.19784232566160803   0.38854653590346255   0.004538366845204598   0.7059017237681704   0.6644651122448769   0.9709065891597194   0.6427941081084465   0.7061839451617736   0.3212763418666171   0.2758188919896954   0.25934804828125796   0.4843552836115978   0.9375812841467397   0.7490776223648652   0.9417036847244622   0.7332492068540001   0.4530438924728307   0.08897629055017457   0.8364067744285404   0.33491481723363425   0.5218485549115143   0.2250680301972847   0.37072757257184547   0.24375748879217607   0.32400622924990624   0.8365214942938222   0.3661892057266409   0.5378557650240057   0.6595411170050293   0.8656149051341027   0.7233950976181944   0.8316718198622322   0.3382647751384122   0.5897960131444073   0.4640470493369364   0.34731653625063436   0.4006834909916725   0.8407183907795421   0.5223433646124742   0.6140673293966342   0.9476395985188418   0.7517421002293675   0.6859365901839338   0.27915251216299997   0.4257910436073275   0.5266740700320829
0.31520901761208836   0.03539502337082389   0.10178481435742125   0.6901525757382607   0.9490198118854475   0.49753925834681817   0.44224369735239194   0.8245376706041581   0.22562471426725306   0.6658674384845861   0.10397892221397975   0.23474165745975079   0.7615776649303166   0.3185509022339517   0.7032954312223073   0.39402326668020865   0.23923430031784237   0.7044835728373174   0.7556558327034655   0.6422811664508411   0.5532977101339086   0.42533106067431753   0.329864789096138   0.11560709641875827   0.23808869252182022   0.38993603730349363   0.22807997473871672   0.42545452068049755   0.28906888063637276   0.8923967789566755   0.7858362773863248   0.6009168500763394   0.0634441663691197   0.2265293404720894   0.681857355172345   0.3661751926165887   0.30186650143880306   0.9079784382381377   0.9785619239500377   0.97215192593638   0.06263220112096068   0.20349486540082024   0.22290609124657226   0.3298707594855389   0.5093344909870522   0.7781638047265027   0.8930413021504343   0.21426366306678063   0.27124579846523195   0.38822776742300913   0.6649613274117175   0.7888091423862831   0.9821769178288592   0.49583098846633367   0.8791250500253929   0.18789229230994361   0.9187327514597394   0.2693016479942443   0.19726769485304785   0.8217170996933549   0.6168662500209364   0.36132320975610654   0.2187057709030101   0.8495651737569749
0.5542340488999757   0.15782834435528634   0.9957996796564379   0.519694414271436   0.04489955791292356   0.3796645396287836   0.10275837750600356   0.30543075120465535   0.7736537594476917   0.9914367722057745   0.43779705009428593   0.5166216088183723   0.7914768416188325   0.4956057837394408   0.5586720000688931   0.3287293165084286   0.872744090159093   0.22630413574519656   0.36140430521584527   0.5070122168150737   0.2558778401381566   0.8649809259890899   0.14269853431283513   0.6574470430580989   0.7016437912381809   0.7071525816338037   0.1468988546563973   0.13775262878666283   0.6567442333252573   0.32748804200502   0.044140477150393743   0.8323218775820075   0.8830904738775658   0.33605126979924554   0.6063434270561078   0.3157002687636352   0.09161363225873326   0.8404454860598047   0.04767142698721467   0.9869709522552066   0.21886954209964024   0.6141413503146081   0.6862671217713694   0.47995873544013284   0.9629917019614835   0.7491604243255182   0.5435685874585342   0.822511692382034   0.26134791072330266   0.042007842691714536   0.39666973280213697   0.6847590635953712   0.6046036773980453   0.7145198006866945   0.3525292556517432   0.8524371860133637   0.7215132035204795   0.378468530887449   0.7461858285956354   0.5367369172497285   0.6298995712617463   0.5380230448276443   0.6985144016084208   0.5497659649945219
0.41103002916210607   0.9238816945130361   0.012247279837051367   0.0698072295543891   0.4480383272006225   0.17472127018751799   0.4686786923785171   0.2472955371723551   0.18669041647731982   0.13271342749580345   0.07200895957638015   0.562536473576984   0.5820867390792746   0.41819362680910893   0.7194797039246369   0.7100992875636203   0.860573535558795   0.039725095921659924   0.9732938753290015   0.17336237031389182   0.2306739642970487   0.5017020510940157   0.2747794737205807   0.6235964053193699   0.8196439351349426   0.5778203565809795   0.26253219388352933   0.5537891757649808   0.3716056079343202   0.4030990863934615   0.7938535015050122   0.3064936385926257   0.18491519145700036   0.2703856588976581   0.7218445419286321   0.7439571650156417   0.6028284523777259   0.8521920320885491   0.002364838003995162   0.03385787745202144   0.7422549168189309   0.8124669361668893   0.02907096267499368   0.8604955071381296   0.5115809525218822   0.3107648850728736   0.754291488954413   0.23689910181875973   0.6919370173869395   0.7329445284918942   0.4917592950708836   0.683109926053779   0.32033140945261934   0.32984544209843264   0.6979057935658713   0.3766162874611533   0.13541621799561898   0.05945978320077456   0.9760612516372393   0.6326591224455115   0.5325877656178931   0.20726775111222542   0.9736964136332441   0.5988012449934901
0.7903328487989624   0.3948008149453362   0.9446254509582505   0.7383057378553605   0.2787518962770802   0.08403592987246258   0.1903339620038375   0.5014066360366007   0.5868148788901407   0.35109140138056844   0.6985746669329539   0.8182967099828218   0.2664834694375214   0.021245959282135823   0.0006688733670824692   0.4416804225216685   0.13106725144190237   0.9617861760813613   0.024607621729843154   0.809021300076157   0.5984794858240092   0.7545184249691359   0.050911208096599   0.21022005508266692   0.8081466370250469   0.35971761002379965   0.10628575713834852   0.4719143172273065   0.5293947407479668   0.2756816801513371   0.9159517951345111   0.9705076811907057   0.942579861857826   0.9245902787707686   0.21737712820155716   0.15221097120788396   0.6760963924203047   0.9033443194886328   0.2167082548344747   0.7105305486862155   0.5450291409784023   0.9415581434072715   0.19210063310463155   0.9015092486100584   0.946549655154393   0.1870397184381357   0.14118942500803253   0.6912891935273915   0.13840301812934616   0.8273221084143361   0.03490366786968401   0.21937487630008506   0.6090082773813794   0.551640428262999   0.11895187273517298   0.24886719510937932   0.6664284155235534   0.6270501494922304   0.9015747445336159   0.09665622390149538   0.9903320231032487   0.7237058300035976   0.6848664896991411   0.38612567521527996
0.4453028821248464   0.7821476865963259   0.4927658565945096   0.48461642660522153   0.4987532269704533   0.5951079681581902   0.35157643158647706   0.79332723307783   0.3603502088411072   0.7677858597438543   0.31667276371679304   0.5739523567777449   0.7513419314597277   0.21614543148085527   0.19772089098162007   0.3250851616683656   0.08491351593617436   0.5890952819886249   0.29614614644800424   0.22842893776687023   0.09458149283292563   0.8653894519850275   0.6112796567488631   0.8423032625515903   0.6492786107080792   0.0832417653887015   0.11851380015435352   0.35768683594636874   0.15052538373762586   0.48813379723051126   0.7669373685678764   0.5643596028685388   0.7901751748965187   0.720347937486657   0.4502646048510834   0.9904072460907938   0.038833243436790926   0.5042025060058017   0.25254371386946334   0.6653220844224282   0.9539197275006166   0.9151072240171767   0.9563975674214591   0.43689314665555795   0.859338234667691   0.04971777203214929   0.34511791067259595   0.5945898841039676   0.21005962395961172   0.9664760066434478   0.22660411051824245   0.2369030481575989   0.059534240221985876   0.47834220941293654   0.459666741950366   0.6725434452890602   0.2693590653254672   0.7579942719262796   0.009402137099282603   0.6821361991982663   0.2305258218886763   0.25379176592047786   0.7568584232298193   0.016814114775838135
0.2766060943880597   0.3386845419033011   0.8004608558083602   0.5799209681202802   0.4172678597203688   0.28896676987115183   0.4553429451357643   0.9853310840163125   0.20720823576075703   0.32249076322770404   0.22873883461752184   0.7484280358587136   0.14767399553877114   0.8441485538147675   0.7690720926671558   0.07588459056965347   0.878314930213304   0.0861542818884879   0.7596699555678732   0.3937483913713871   0.6477891083246277   0.83236251596801   0.0028115323380539558   0.376934276595549   0.37118301393656794   0.4936779740647089   0.20235067652969374   0.7970133084752689   0.9539151542161992   0.20471120419355712   0.7470077313939294   0.8116822244589563   0.7467069184554421   0.8822204409658531   0.5182688967764076   0.06325418860024269   0.599032922916671   0.03807188715108566   0.7491968041092517   0.9873695980305892   0.7207179927033671   0.9519176052625977   0.9895268485413785   0.593621206659202   0.07292888437873941   0.11955508929458773   0.9867153162033245   0.21668693006365308   0.7017458704421715   0.6258771152298788   0.7843646396736308   0.4196736215883843   0.7478307162259723   0.42116591103632167   0.03735690827970138   0.607991397129428   0.0011237977705301355   0.5389454700704686   0.5190880115032938   0.5447372085291853   0.40209087485385914   0.5008735829193829   0.769891207394042   0.5573676104985961
0.6813728821504921   0.5489559776567852   0.7803643588526635   0.9637464038393939   0.6084439977717526   0.4294008883621974   0.7936490426493389   0.7470594737757409   0.9066981273295812   0.8035237731323186   0.009284402975708098   0.3273858521873566   0.15886741110360889   0.382357862095997   0.9719274946960067   0.7193944550579287   0.15774361333307874   0.8434123920255284   0.45283948319271294   0.17465724652874337   0.7556527384792197   0.3425388091061455   0.6829482757986709   0.6172896360301473   0.07427985632872756   0.7935828314493604   0.9025839169460075   0.6535432321907534   0.4658358585569749   0.36418194308716295   0.10893487429666852   0.9064837584150125   0.5591377312273937   0.5606581699548443   0.09965047132096043   0.5790979062276559   0.4002703201237849   0.17830030785884735   0.12772297662495372   0.8597034511697272   0.24252670679070612   0.33488791583331895   0.6748834934322407   0.6850462046409839   0.4868739683114865   0.9923491067271735   0.9919352176335698   0.06775656861083654   0.41259411198275897   0.19876627527781313   0.08935130068756236   0.4142133364200832   0.946758253425784   0.8345843321906502   0.9804164263908939   0.5077295780050707   0.38762052219839027   0.27392616223580585   0.8807659550699334   0.9286316717774147   0.9873502020746054   0.09562585437695852   0.7530429784449797   0.06892822060768745
0.7448234952838992   0.7607379385436396   0.07815948501273894   0.38388201596670357   0.2579495269724128   0.7683888318164661   0.08622426737916913   0.316125447355867   0.8453554149896538   0.569622556538653   0.9968729666916067   0.9019121109357838   0.8985971615638698   0.7350382243480028   0.01645654030071294   0.39418253293071326   0.5109766393654795   0.4611120621121969   0.13569058523077954   0.4655508611532985   0.5236264372908741   0.3654862077352384   0.38264760678579984   0.3966226405456111   0.7788029420069749   0.6047482691915989   0.3044881217730609   0.0127406245789075   0.5208534150345621   0.8363594373751327   0.21826385439389176   0.6966151772230404   0.6754980000449082   0.2667368808364798   0.221390887702285   0.7947030662872566   0.7769008384810384   0.531698656488477   0.20493434740157207   0.40052053335654336   0.26592419911555887   0.0705865943762801   0.06924376217079252   0.9349696722032449   0.7422977618246848   0.7051003866410417   0.6865961553849926   0.5383470316576338   0.9634948198177099   0.10035211744944286   0.3821080336119318   0.5256064070787263   0.4426414047831479   0.2639926800743101   0.16384417921804   0.8289912298556859   0.7671434047382397   0.9972557992378303   0.942453291515755   0.03428816356842921   0.9902425662572013   0.4655571427493533   0.737518944114183   0.6337676302118859
0.7243183671416424   0.39497054837307316   0.6682751819433904   0.698797958008641   0.9820206053169577   0.6898701617320314   0.9816790265583978   0.16045092635100713   0.01852578549924769   0.5895180442825886   0.599570992946466   0.6348445192722808   0.5758843807160998   0.3255253642082785   0.435726813728426   0.8058532894165951   0.8087409759778601   0.3282695649704482   0.49327352221267096   0.7715651258481658   0.8184984097206588   0.8627124222210949   0.755754578098488   0.13779749563627997   0.09418004257901637   0.46774187384802174   0.08747939615509755   0.43899953762763905   0.11215943726205872   0.7778717121159903   0.10580036959669979   0.2785486112766319   0.09363365176281103   0.18835366783340166   0.5062293766502338   0.6437040920043511   0.5177492710467112   0.8628283036251232   0.07050256292180787   0.837850802587756   0.7090082950688512   0.534558738654675   0.5772290407091369   0.06628567673959022   0.8905098853481924   0.6718463164335801   0.8214744626106489   0.9284881811033102   0.7963298427691761   0.20410444258555832   0.7339950664555513   0.4894886434756712   0.6841704055071173   0.42623273046956806   0.6281946968588517   0.21094003219903937   0.5905367537443063   0.2378790626361664   0.12196532020861778   0.5672359401946884   0.07278748269759502   0.37505075901104323   0.051462757286809914   0.7293851376069322
0.36377918762874384   0.8404920203563683   0.474233716577673   0.6630994608673421   0.4732693022805515   0.16864570392278821   0.6527592539670241   0.7346112797640318   0.6769394595113755   0.9645412613372298   0.9187641875114726   0.24512263628836056   0.9927690540042581   0.5383085308676618   0.29056949065262105   0.03418260408932121   0.4022323002599518   0.3004294682314954   0.16860417044400328   0.4669466638946329   0.32944481756235683   0.9253787092204522   0.11714141315719336   0.7375615262877006   0.9656656299336129   0.0848866888640839   0.6429076965795204   0.07446206542035853   0.4923963276530615   0.9162409849412957   0.9901484426124963   0.33985078565632676   0.815456868141686   0.9516997236040659   0.07138425510102366   0.09472814936796617   0.822687814137428   0.413391192736404   0.7808147644484026   0.060545545278644954   0.4204555138774761   0.11296172450490859   0.6122105940043994   0.5935988813840121   0.09101069631511928   0.18758301528445642   0.495069180847206   0.8560373550963115   0.1253450663815063   0.1026963264203725   0.8521614842676857   0.7815752896759529   0.6329487387284448   0.1864553414790768   0.8620130416551893   0.4417245040196262   0.8174918705867587   0.234755617875011   0.7906287865541657   0.34699635465166   0.9948040564493308   0.821364425138607   0.009814022105763051   0.2864508093730151
0.5743485425718546   0.7084027006336985   0.3976034281013637   0.692851927989003   0.48333784625673537   0.5208196853492421   0.9025342472541577   0.8368145728926916   0.35799277987522904   0.41812335892886954   0.050372762986472065   0.055239283216738606   0.7250440411467842   0.2316680174497927   0.18835972133128273   0.6135147791971124   0.9075521705600256   0.9969123995747817   0.3977309347771171   0.2665184245454524   0.9127481141106948   0.17554797443617468   0.38791691267135403   0.9800676151724372   0.33839957153884015   0.4671452738024763   0.9903134845699904   0.28721568718343427   0.8550617252821048   0.9463255884532342   0.08777923731583262   0.45040111429074275   0.4970689454068758   0.5282022295243647   0.03740647432936055   0.39516183107400416   0.7720249042600915   0.29653421207457203   0.8490467529980779   0.7816470518768918   0.8644727337000659   0.29962181249979036   0.45131581822096073   0.5151286273314394   0.9517246195893712   0.12407383806361566   0.06339890554960671   0.535061012159002   0.613325048050531   0.6569285642611394   0.0730854209796164   0.2478453249755678   0.7582633227684261   0.7106029758079052   0.9853061836637838   0.7974442106848251   0.2611943773615504   0.18240074628354044   0.9478997093344232   0.4022823796108209   0.48916947310145886   0.8858665342089684   0.09885295633634543   0.6206353277339292
0.6246967394013929   0.5862447217091781   0.6475371381153847   0.10550670040248984   0.6729721198120218   0.4621708836455624   0.584138232565778   0.5704456882434877   0.05964707176149082   0.805242319384423   0.5110528115861616   0.32260036326791997   0.3013837489930647   0.09463934357651786   0.5257466279223778   0.5251561525830949   0.0401893716315143   0.9122385972929774   0.5778469185879546   0.122873772972274   0.5510198985300554   0.026372063084009   0.4789939622516091   0.5022384452383448   0.9263231591286625   0.4401273413748309   0.8314568241362245   0.396731744835855   0.2533510393166407   0.9779564577292685   0.24731859157044647   0.8262860565923672   0.1937039675551499   0.17271413834484547   0.7362657799842849   0.5036856933244472   0.8923202185620852   0.07807479476832761   0.21051915206190713   0.9785295407413523   0.852130846930571   0.1658361974753502   0.6326722334739525   0.8556557677690783   0.3011109484005155   0.1394641343913412   0.15367827122234343   0.3534173225307335   0.37478778927185297   0.6993367930165103   0.322221447086119   0.9566855776948785   0.12143674995521225   0.7213803352872418   0.07490285551567252   0.13039952110251132   0.9277327824000623   0.5486661969423963   0.3386370755313876   0.6267138277780641   0.0354125638379771   0.4705914021740687   0.12811792346948048   0.6481842870367118
0.18328171690740616   0.30475520469871853   0.4954456899955279   0.7925285192676335   0.8821707685068907   0.1652910703073773   0.3417674187731845   0.43911119673689997   0.5073829792350377   0.465954277290867   0.01954597168706549   0.48242561904202147   0.38594622927982547   0.7445739420036253   0.944643116171393   0.3520260979395101   0.4582134468797631   0.1959077450612289   0.6060060406400054   0.7253122701614461   0.422800883041786   0.7253163428871602   0.4778881171705249   0.07712798312473425   0.23951916613437985   0.4205611381884417   0.982442427174997   0.2845994638571008   0.35734839762748916   0.2552700678810644   0.6406750084018125   0.8454882671202008   0.8499654183924514   0.7893157905901974   0.621129036714747   0.36306264807817934   0.464019189112626   0.04474184858657215   0.676485920543354   0.011036550138669225   0.005805742232862918   0.8488341035253433   0.07047987990334864   0.2857242799772232   0.5830048591910769   0.12351776063818305   0.5925917627328238   0.20859629685248895   0.3434856930566971   0.7029566224497413   0.6101493355578268   0.9239968329953882   0.9861372954292079   0.44768655456867695   0.9694743271560143   0.07850856587518738   0.13617187703675646   0.6583707639784796   0.3483452904412674   0.7154459177970081   0.6721526879241304   0.6136289153919074   0.6718593698979134   0.7044093676583388
0.6663469456912675   0.7647948118665642   0.6013794899945647   0.4186850876811156   0.08334208650019059   0.6412770512283811   0.008787727261740944   0.21008879082862666   0.7398563934434935   0.9383204287786397   0.39863839170391413   0.2860919578332385   0.7537190980142856   0.4906338742099628   0.4291640645478998   0.2075833919580511   0.6175472209775291   0.8322631102314832   0.08081877410663243   0.4921374741610431   0.9453945330533987   0.2186341948395758   0.40895940420871907   0.7877281065027042   0.2790475873621312   0.45383938297301163   0.8075799142141544   0.36904301882158863   0.19570550086194063   0.8125623317446306   0.7987921869524134   0.15895422799296197   0.45584910741844714   0.8742419029659907   0.4001537952484993   0.8728622701597235   0.7021300094041615   0.38360802875602795   0.9709897307005995   0.6652788782016723   0.08458278842663237   0.5513449185245447   0.890170956593967   0.1731414040406293   0.13918825537323365   0.3327107236849689   0.481211552385248   0.3854132975379251   0.8601406680111024   0.8788713407119573   0.6736316381710936   0.016370278716336433   0.6644351671491618   0.06630900896732678   0.8748394512186801   0.8574160507233745   0.20858605973071467   0.19206710600133603   0.47468565597018086   0.9845537805636511   0.5064560503265532   0.8084590772453081   0.5036959252695814   0.31927490236197864
0.4218732618999208   0.2571141587207634   0.6135249686756143   0.14613349832134934   0.28268500652668715   0.9244034350357945   0.13231341629036633   0.7607202007834243   0.4225443385155847   0.045532094323837174   0.45868177811927274   0.7443499220670878   0.7581091713664229   0.9792230853565104   0.5838423269005926   0.8869338713437134   0.5495231116357082   0.7871559793551743   0.10915667093041168   0.9023800907800623   0.04306706130915507   0.9786969021098663   0.6054607456608303   0.5831051884180837   0.6211937994092342   0.7215827433891029   0.991935776985216   0.43697169009673437   0.33850879288254715   0.7971793083533085   0.8596223606948497   0.67625148931331   0.9159644543669625   0.7516472140294713   0.4009405825755769   0.9319015672462222   0.15785528300053955   0.7724241286729608   0.8170982556749844   0.044967695902508834   0.6083321713648313   0.9852681493177865   0.7079415847445727   0.14258760512244648   0.5652651100556763   0.006571247207920211   0.1024808390837424   0.5594824167043627   0.944071310646442   0.2849885038188173   0.11054506209852642   0.12251072660762838   0.6055625177638948   0.4878091954655088   0.2509227014036768   0.4462592372943183   0.6895980633969323   0.7361619814360375   0.8499821188280998   0.5143576700480961   0.5317427803963928   0.9637378527630767   0.03288386315311547   0.46938997414558725
0.9234106090315615   0.9784697034452902   0.3249422784085428   0.3268023690231408   0.35814549897588516   0.9718984562373699   0.22246143932480036   0.767319952318778   0.4140741883294432   0.6869099524185526   0.11191637722627393   0.6448092257111496   0.8085116705655484   0.1991007569530438   0.8609936758225971   0.19854998841683136   0.11891360716861604   0.4629387755170063   0.011011556994497313   0.6841923183687353   0.5871708267722233   0.4992009227539297   0.9781276938413819   0.214802344223148   0.6637602177406619   0.5207312193086395   0.653185415432839   0.8879999752000072   0.30561471876477664   0.5488327630712696   0.4307239761080387   0.12068002288122916   0.8915405304353334   0.861922810652717   0.3188075988817648   0.47587079717007946   0.08302885986978506   0.6628220536996732   0.4578139230591676   0.2773208087532481   0.964115252701169   0.1998832781826669   0.44680236606467033   0.5931284903845129   0.3769444259289457   0.7006823554287372   0.46867467222328846   0.37832614616136484   0.7131842081882839   0.1799511361200977   0.8154892567904494   0.4903261709613576   0.40756948942350724   0.631118373048828   0.38476528068241067   0.36964614808012847   0.5160289589881738   0.7691955623961111   0.06595768180064589   0.893775350910049   0.43300009911838877   0.10637350869643784   0.6081437587414783   0.6164545421568008
0.4688848464172197   0.906490230513771   0.16134139267680794   0.023326051772288046   0.09194042048827399   0.20580787508503373   0.6926667204535194   0.6449999056109232   0.37875621229999007   0.025856738964936038   0.87717746366307   0.15467373464956558   0.9711867228764828   0.394738365916108   0.49241218298065936   0.785027586569437   0.455157763888309   0.6255428035199969   0.4264545011800135   0.891252235659388   0.022157664769920257   0.5191692948235591   0.8183107424385352   0.2747976935025872   0.5532728183527005   0.6126790643097881   0.6569693497617273   0.2514716417302991   0.46133239786442654   0.4068711892247544   0.9643026293082079   0.6064717361193759   0.08257618556443647   0.3810144502598184   0.0871251656451378   0.45179800146981036   0.11138946268795366   0.9862760843437104   0.5947129826644785   0.6667704149003733   0.6562316987996447   0.3607332808237135   0.16825848148446493   0.7755181792409852   0.6340740340297244   0.8415639860001544   0.3499477390459297   0.500720485738398   0.08080121567702388   0.22888492169036623   0.6929783892842024   0.24924884400809885   0.6194688178125973   0.8220137324656118   0.7286757599759945   0.6427771078887229   0.5368926322481609   0.44099928220579343   0.6415505943308567   0.19097910641891255   0.42550316956020723   0.45472319786208304   0.046837611666378315   0.5242086915185393
0.7692714707605626   0.09398991703836956   0.8785791301819134   0.7486905122775541   0.13519743673083814   0.2524259310382152   0.5286313911359837   0.2479700265391561   0.05439622105381427   0.023541009347848994   0.8356530018517813   0.9987211825310572   0.4349274032412169   0.2015272768822372   0.10697724187578674   0.3559440746423343   0.8980347709930561   0.7605279946764438   0.46542664754493   0.16496496822342174   0.47253160143284884   0.3058047968143608   0.4185890358785517   0.6407562767048824   0.7032601306722863   0.2118148797759912   0.5400099056966383   0.8920657644273283   0.5680626939414481   0.959388948737776   0.011378514560654616   0.6440957378881723   0.5136664728876339   0.935847939389927   0.17572551270887335   0.6453745553571151   0.07873906964641697   0.7343206625076898   0.0687482708330866   0.2894304807147807   0.1807042986533609   0.973792667831246   0.6033216232881566   0.12446551249135898   0.708172697220512   0.6679878710168853   0.18473258740960494   0.4837092357864765   0.004912566548225768   0.45617299124089405   0.6447226817129666   0.5916434713591482   0.4368498726067776   0.49678404250311803   0.633344167152312   0.9475477334709759   0.9231833997191438   0.560936103113191   0.4576186544434387   0.3021731781138608   0.8444443300727268   0.8266154406055012   0.3888703836103521   0.012742697399080084
0.6637400314193659   0.8528227727742552   0.7855487603221954   0.8882771849077211   0.9555673341988538   0.18483490175737   0.6008161729125906   0.4045679491212446   0.9506547676506281   0.728661910516476   0.956093491199624   0.8129244777620964   0.5138048950438504   0.2318778680133579   0.3227493240473119   0.8653767442911205   0.5906214953247066   0.6709417649001669   0.8651306696038732   0.5632035661772598   0.74617716525198   0.8443263242946657   0.4762602859935211   0.5504608687781797   0.08243713383261407   0.9915035515204105   0.6907115256713257   0.6621836838704586   0.1268697996337603   0.8066686497630404   0.08989535275873507   0.257615734749214   0.1762150319831323   0.0780067392465645   0.13380186155911117   0.44469125698711753   0.6624101369392819   0.8461288712332066   0.8110525375117993   0.579314512695997   0.07178864161457521   0.1751871063330397   0.9459218679079261   0.016110946518737176   0.3256114763625953   0.330860782038374   0.46966158191440505   0.4656500777405575   0.2431743425299812   0.33935723051796357   0.7789500562430794   0.8034663938700989   0.11630454289622093   0.5326885807549231   0.6890547034843444   0.5458506591208849   0.9400895109130887   0.4546818415083586   0.5552528419252332   0.10115940213376735   0.27767937397380676   0.6085529702751521   0.7442003044134339   0.5218448894377704
0.20589073235923155   0.4333658639421124   0.7982784365055078   0.5057339429190332   0.8802792559966363   0.10250508190373837   0.3286168545911027   0.040083865178475744   0.6371049134666551   0.7631478513857748   0.5496667983480233   0.23661747130837685   0.5208003705704342   0.23045927063085167   0.860612094863679   0.6907668121874919   0.5807108596573455   0.775777429122493   0.3053592529384458   0.5896074100537246   0.3030314856835387   0.16722445884734097   0.5611589485250119   0.06776252061595418   0.09714075332430715   0.7338585949052285   0.7628805120195042   0.5620285776969209   0.21686149732767088   0.6313535130014902   0.4342636574284015   0.5219447125184452   0.5797565838610158   0.8682056616157154   0.8845968590803782   0.28532724121006836   0.05895621329058172   0.6377463909848637   0.02398476421669926   0.5945604290225764   0.4782453536332362   0.8619689618623707   0.7186255112782535   0.004953018968851829   0.17521386794969754   0.6947445030150298   0.1574665627532415   0.9371904983528977   0.07807311462539038   0.9608859081098011   0.3945860507337373   0.3751619206559767   0.8612116172977196   0.32953239510831095   0.9603223933053358   0.8532172081375314   0.28145503343670364   0.4613267334925955   0.07572553422495756   0.5678899669274631   0.22249882014612196   0.8235803425077318   0.051740770008258295   0.9733295379048867
0.7442534665128857   0.9616113806453611   0.33311525873000486   0.9683765189360348   0.5690395985631882   0.2668668776303313   0.17564869597676333   0.03118602058313723   0.4909664839377978   0.30598096952053017   0.781062645243026   0.6560240999271605   0.6297548666400783   0.9764485744122192   0.8207402519376903   0.802806891789629   0.3482998332033746   0.5151218409196237   0.7450147177127326   0.23491692486216592   0.12580101305725266   0.6915414984118919   0.6932739477044744   0.26158738695727923   0.38154754654436696   0.7299301177665308   0.36015868897446957   0.29321086802124435   0.8125079479811788   0.46306324013619954   0.18450999299770623   0.2620248474381071   0.321541464043381   0.15708227061566937   0.4034473477546802   0.6060007475109466   0.6917865974033027   0.18063369620345016   0.58270709581699   0.8031938557213175   0.34348676419992813   0.6655118552838265   0.8376923781042572   0.5682769308591515   0.21768575114267544   0.9739703568719346   0.14441843039978286   0.30668954390187236   0.8361382045983085   0.24404023910540373   0.7842597414253133   0.013478675880628031   0.02363025661712967   0.7809769989692043   0.5997497484276071   0.751453828442521   0.7020887925737487   0.6238947283535349   0.19630240067292687   0.14545308093157433   0.010302195170445932   0.44326103215008467   0.6135953048559369   0.3422592252102568
0.6668154309705179   0.7777491768662582   0.7759029267516797   0.7739822943511052   0.4491296798278424   0.8037788199943237   0.6314844963518969   0.46729275044923285   0.6129914752295339   0.5597385808889199   0.8472247549265836   0.4538140745686048   0.5893612186124042   0.7787615819197157   0.24747500649897647   0.7023602461260839   0.8872724260386556   0.15486685356618085   0.051172605826049586   0.5569071651945096   0.8769702308682097   0.7116058214160962   0.43757730097011266   0.21464793998425274   0.21015479989769184   0.933856644549838   0.661674374218433   0.44066564563314753   0.7610251200698495   0.1300778245555144   0.030189877866536152   0.9733728951839147   0.14803364484031553   0.5703392436665945   0.18296512293995262   0.5195588206153099   0.5586724262279112   0.7915776617468788   0.9354901164409761   0.817198574489226   0.6714000001892557   0.636710808180698   0.8843175106149266   0.2602914092947164   0.794429769321046   0.9251049867646018   0.4467402096448139   0.045643469310463675   0.5842749694233541   0.9912483422147639   0.785065835426381   0.6049778236773161   0.8232498493535048   0.8611705176592495   0.7548759575598448   0.6316049284934014   0.6752162045131892   0.2908312739926549   0.5719108346198921   0.1120461078780916   0.11654377828527793   0.4992536122457761   0.636420718178916   0.29484753338886566
0.4451437780960223   0.8625428040650781   0.7521032075639894   0.034556124094149224   0.6507140087749763   0.9374378173004763   0.3053629979191755   0.9889126547836855   0.06643903935162211   0.9461894750857124   0.5202971624927946   0.3839348311063694   0.2431891899981174   0.08501895742646297   0.7654212049329497   0.752329902612968   0.5679729854849282   0.7941876834338081   0.1935103703130576   0.6402837947348763   0.4514292071996503   0.29493407118803194   0.5570896521341416   0.3454362613460107   0.006285429103628007   0.4323912671229539   0.8049864445701521   0.3108801372518615   0.35557142032865174   0.49495344982247763   0.49962344665097663   0.3219674824681759   0.28913238097702965   0.5487639747367652   0.9793262841581821   0.9380326513618065   0.04594319097891224   0.46374501731030227   0.21390507922523233   0.18570274874883858   0.47797020549398406   0.6695573338764942   0.020394708912174743   0.5454189540139622   0.026540998294333765   0.37462326268846224   0.46330505677803313   0.19998269266795157   0.020255569190705758   0.9422319955655084   0.658318612207881   0.8891025554160901   0.6646841488620541   0.4472785457430307   0.15869516555690433   0.5671350729479142   0.37555176788502437   0.8985145710062655   0.17936888139872223   0.6291024215861077   0.32960857690611217   0.43476955369596326   0.9654638021734899   0.4433996728372691
0.8516383714121281   0.7652122198194691   0.9450690932613152   0.8979807188233069   0.8250973731177943   0.3905889571310068   0.48176403648328203   0.6979980261553553   0.8048418039270886   0.44835696156549837   0.823445424275401   0.8088954707392652   0.14015765506503455   0.0010784158224676488   0.6647502587184967   0.24176039779135097   0.7646058871800102   0.10256384481620212   0.48538137731977443   0.6126579762052433   0.43499731027389804   0.6677942911202389   0.5199175751462846   0.16925830336797418   0.5833589388617699   0.9025820713007698   0.5748484818849694   0.2712775845446673   0.7582615657439756   0.511993114169763   0.09308444540168735   0.573279558389312   0.953419761816887   0.06363615260426465   0.26963902112628635   0.7643840876500468   0.8132621067518524   0.062557736781797   0.6048887624077897   0.5226236898586958   0.04865621957184225   0.9599938919655949   0.11950738508801524   0.9099657136534526   0.6136589092979442   0.292199600845356   0.5995898099417307   0.7407074102854784   0.03029997043617429   0.38961752954458617   0.024741328056761363   0.46942982574081105   0.2720384046921987   0.8776244153748232   0.9316568826550741   0.896150267351499   0.3186186428753117   0.8139882627705585   0.6620178615287877   0.13176617970145224   0.5053565361234593   0.7514305259887615   0.057129099120998006   0.6091424898427564
0.456700316551617   0.7914366340231667   0.9376217140329828   0.6991767761893039   0.8430414072536728   0.4992370331778106   0.33803190409125206   0.9584693659038255   0.8127414368174986   0.10961950363322441   0.3132905760344907   0.48903954016301443   0.5407030321252998   0.23199508825840126   0.38163369337941666   0.5928892728115154   0.2220843892499881   0.4180068254878428   0.7196158318506289   0.4611230931100631   0.7167278531265289   0.6665762994990813   0.662486732729631   0.8519806032673067   0.2600275365749118   0.8751396654759147   0.7248650186966482   0.15280382707800286   0.416986129321239   0.3759026322981041   0.38683311460539616   0.19433446117417738   0.6042446925037405   0.2662831286648797   0.07354253857090548   0.705294921011163   0.06354166037844067   0.0342880404064784   0.6919088451914888   0.11240564819964764   0.8414572711284526   0.6162812149186356   0.9722930133408598   0.6512825550895845   0.12472941800192373   0.9497049154195543   0.30980628061122883   0.7993019518222778   0.8647018814270119   0.07456524994363962   0.5849412619145806   0.6464981247442749   0.4477157521057729   0.6986626176455355   0.19810814730918447   0.4521636635700976   0.8434710596020324   0.43237948898065587   0.12456560873827897   0.7468687425589345   0.7799293992235917   0.39809144857417744   0.43265676354679017   0.6344630943592869
0.9384721280951392   0.7818102336555418   0.46036375020593034   0.9831805392697024   0.8137427100932155   0.8321053182359875   0.1505574695947015   0.18387858744742458   0.9490408286662035   0.7575400682923479   0.5656162076801209   0.5373804627031497   0.5013250765604307   0.05887745064681237   0.3675080603709364   0.08521679913305205   0.6578540169583982   0.6264979616661566   0.24294245163265746   0.3383480565741175   0.8779246177348065   0.22840651309197904   0.8102856880858673   0.7038849622148305   0.9394524896396672   0.4465962794364372   0.349921937879937   0.7207044229451282   0.12570977954645174   0.6144909612004497   0.19936446828523544   0.5368258354977036   0.17666895088024817   0.8569508929081018   0.6337482606051146   0.999445372794554   0.6753438743198176   0.7980734422612894   0.2662402002341781   0.9142285736615019   0.017489857361419312   0.1715754805951329   0.023297748601520646   0.5758805170873844   0.13956523962661288   0.9431689675031538   0.21301206051565336   0.8719955548725539   0.20011274998694567   0.4965726880667166   0.8630901226357164   0.15129113192742574   0.07440297044049393   0.882081726866267   0.6637256543504809   0.6144652964297221   0.8977340195602458   0.02513083395816517   0.029977393745366402   0.6150199236351681   0.22239014524042824   0.22705739169687578   0.7637371935111883   0.7007913499736662
0.20490028787900894   0.055481911101742894   0.7404394449096676   0.12491083288628174   0.06533504825239606   0.11231294359858907   0.5274273843940143   0.2529152780137279   0.8652222982654504   0.6157402555318724   0.6643372617582979   0.10162414608630212   0.7908193278249565   0.7336585286656055   0.0006116074078169522   0.48715884965657996   0.8930853082647107   0.7085276947074404   0.9706342136624505   0.8721389260214119   0.6706951630242824   0.48147030301056454   0.20689702015126227   0.17134757604774564   0.4657948751452735   0.42598839190882165   0.4664575752415946   0.046436743161463886   0.40045982689287746   0.3136754483102326   0.9390301908475803   0.793521465147736   0.535237528627427   0.6979351927783601   0.27469292908928244   0.6918973190614339   0.7444182008024706   0.9642766641127547   0.2740813216814655   0.20473846940485393   0.8513328925377599   0.25574896940531433   0.3034471080190149   0.3325995433834421   0.18063772951347745   0.7742786663947497   0.09655008786775265   0.16125196733569647   0.7148428543682039   0.3482902744859281   0.6300925126261581   0.1148152241742326   0.31438302747532654   0.0346148261756955   0.6910623217785777   0.32129375902649654   0.7791454988478995   0.33667963339733536   0.4163693926892953   0.6293964399650627   0.03472729804542889   0.3724029692845807   0.14228807100782984   0.4246579705602087
0.183394405507669   0.11665399987926638   0.8388409629888149   0.09205842717676657   0.0027566759941915334   0.3423753334845166   0.7422908751210623   0.9308064598410701   0.28791382162598755   0.9940850589985886   0.11219836249490422   0.8159912356668375   0.973530794150661   0.959470232822893   0.4211360407163265   0.49469747664034097   0.19438529530276158   0.6227905994255577   0.004766648027031212   0.8653010366752784   0.15965799725733268   0.250387630140977   0.8624785770192014   0.44064306611506965   0.9762635917496637   0.1337336302617106   0.02363761403038647   0.34858463893830305   0.9735069157554722   0.7913582967771939   0.2813467389093242   0.41777817909723297   0.6855930941294845   0.7972732377786055   0.16914837641442   0.6017869434303955   0.7120622999788235   0.8378030049557125   0.7480123356980934   0.1070894667900545   0.5176770046760619   0.21501240553015477   0.7432456876710622   0.2417884301147762   0.3580190074187293   0.9646247753891778   0.8807671106518609   0.8011453639997066   0.38175541566906557   0.8308911451274672   0.8571294966214744   0.4525607250614035   0.4082484999135934   0.039532848350273216   0.5757827577121502   0.034782545964170505   0.7226554057841088   0.24225961057166776   0.4066343812977302   0.43299560253377506   0.010593105805285288   0.4044566056159553   0.6586220455996368   0.3259061357437205
0.49291610112922335   0.18944420008580054   0.9153763579285745   0.08411770562894436   0.13489709371049405   0.22481942469662275   0.034609247276713585   0.2829723416292378   0.7531416780414285   0.39392827956915555   0.17747975065523916   0.8304116165678344   0.34489317812783504   0.35439543121888234   0.601696992943089   0.7956290706036638   0.6222377723437262   0.11213582064721458   0.19506261164535876   0.3626334680698888   0.611644666538441   0.7076792150312593   0.536440566045722   0.036727332326168254   0.11872856540921761   0.5182350149454588   0.6210642081171476   0.9526096266972239   0.9838314716987235   0.29341559024883596   0.5864549608404339   0.6696372850679861   0.23068979365729508   0.8994873106796805   0.4089752101851948   0.8392256685001518   0.88579661552946   0.5450918794607981   0.8072782172421058   0.043596597896487926   0.2635588431857338   0.4329560588135835   0.612215605596747   0.6809631298265991   0.6519141766472929   0.7252768437823243   0.07577503955102505   0.6442357975004309   0.5331856112380752   0.20704182883686553   0.4547108314338775   0.691626170803207   0.5493541395393516   0.9136262385880296   0.8682558705934436   0.02198888573522089   0.31866434588205655   0.014138927908349122   0.4592806604082488   0.18276321723506914   0.43286773035259657   0.469047048447551   0.652002443166143   0.1391666193385812
0.16930888716686276   0.036090989633967514   0.03978683756939587   0.4582034895119821   0.5173947105195699   0.31081414585164324   0.9640117980183708   0.8139676920115512   0.9842090992814947   0.10377231701477774   0.5093009665844933   0.12234152120834418   0.434854959742143   0.1901460784267482   0.6410450959910498   0.1003526354731233   0.11619061386008644   0.17600715051839907   0.181764435582801   0.9175894182380542   0.6833228835074899   0.706960102070848   0.5297619924166581   0.778422798899473   0.5140139963406272   0.6708691124368805   0.48997515484726223   0.3202193093874909   0.9966192858210572   0.3600549665852373   0.5259633568288914   0.5062516173759397   0.01241018653956251   0.25628264957045954   0.01666239024439807   0.3839100961675955   0.5775552267974194   0.06613657114371133   0.3756172942533483   0.28355746069447224   0.46136461293733305   0.8901294206253123   0.1938528586705473   0.36596804245641806   0.7780417294298432   0.18316931855446422   0.6640908662538892   0.5875452435569452   0.264027733089216   0.5123002061175838   0.17411571140662702   0.2673259341694542   0.2674084472681588   0.15224523953234645   0.6481523545777357   0.7610743167935144   0.2549982607285963   0.8959625899618869   0.6314899643333376   0.377164220625919   0.6774430339311769   0.8298260188181756   0.25587267007998926   0.09360675993144674
0.2160784209938438   0.9396965981928633   0.06201981140944197   0.7276387174750286   0.43803669156400066   0.756527279638399   0.39792894515555277   0.14009347391808355   0.17400895847478462   0.24422707352081538   0.22381323374892573   0.8727675397486293   0.9066005112066258   0.09198183398846894   0.5756608791711901   0.11169322295511486   0.6516022504780294   0.196019244026582   0.9441709148378525   0.7345290023291959   0.9741592165468527   0.3661932252084064   0.6882982447578633   0.6409222423977492   0.7580807955530088   0.4264966270155431   0.6262784333484213   0.9132835249227205   0.3200441039890082   0.669969347377144   0.22834948819286854   0.7731900510046369   0.14603514551422359   0.42574227385632857   0.004536254443942812   0.9004225112560076   0.2394346343075978   0.33376043986785964   0.4288753752727527   0.7887292883008927   0.5878323838295684   0.13774119584127764   0.48470446043490023   0.05420028597169683   0.6136731672827157   0.7715479706328713   0.796406215677037   0.41327804357394765   0.8555923717297069   0.34505134361732814   0.17012778232861567   0.4999945186512272   0.5355482677406987   0.6750819962401842   0.9417782941357471   0.7268044676465902   0.38951312222647516   0.24933972238385563   0.9372420396918043   0.8263819563905827   0.15007848791887735   0.915579282515996   0.5083666644190517   0.037652668089689936
0.562246104089309   0.7778380866747183   0.02366220398415139   0.9834523821179931   0.9485729368065933   0.006290116041847118   0.22725598830711444   0.5701743385440454   0.09298056507688636   0.661238772424519   0.057128205978498756   0.07017981989281827   0.5574322973361876   0.9861567761843347   0.11534991184275162   0.343375352246228   0.1679191751097125   0.7368170538004791   0.17810787215094728   0.5169933958556454   0.01784068719083513   0.8212377712844832   0.6697412077318957   0.47934072776595543   0.4555945831015261   0.04339968460976483   0.6460790037477443   0.49588834564796236   0.5070216462949328   0.037109568567917715   0.4188230154406299   0.9257140071039169   0.4140410812180465   0.37587079614339874   0.3616948094621311   0.8555341872110986   0.8566087838818589   0.38971401995906396   0.2463448976193795   0.5121588349648706   0.6886896087721464   0.6528969661585848   0.0682370254684322   0.9951654391092252   0.6708489215813113   0.8316591948741017   0.39849581773653653   0.5158247113432698   0.21525433847978512   0.7882595102643368   0.7524168139887922   0.01993636569530744   0.7082326921848523   0.7511499416964191   0.33359379854816235   0.09422235859139055   0.29419161096680574   0.37527914555302033   0.9718989890860312   0.2386881713802919   0.4375828270849469   0.9855651255939564   0.7255540914666517   0.7265293364154213
0.7488932183128005   0.33266815943537154   0.6573170659982196   0.7313638973061961   0.07804429673148924   0.5010089645612699   0.258821248261683   0.21553918596292634   0.8627899582517041   0.712749454296933   0.5064044342728908   0.1956028202676189   0.15455726606685186   0.9615995126005139   0.17281063572472846   0.10138046167622836   0.860365655100046   0.5863203670474936   0.2009116466386972   0.8626922902959364   0.4227828280150992   0.6007552414535372   0.4753575551720455   0.1361629538805151   0.6738896097022987   0.2680870820181657   0.8180404891738259   0.40479905657431897   0.5958453129708094   0.7670781174568958   0.5592192409121429   0.18925987061139266   0.7330553547191053   0.05432866315996278   0.052814806639252074   0.9936570503437737   0.5784980886522535   0.09272915055944882   0.8800041709145237   0.8922765886675454   0.7181324335522073   0.5064087835119552   0.6790925242758264   0.029584298371608968   0.2953496055371082   0.905653542058418   0.20373496910378094   0.8934213444910939   0.6214599958348095   0.6375664600402522   0.38569447992995504   0.48862228791677487   0.025614682864000055   0.8704883425833564   0.8264752390178122   0.29936241730538227   0.2925593281448947   0.8161596794233936   0.7736604323785601   0.3057053669616085   0.7140612394926412   0.7234305288639448   0.8936562614640364   0.4134287782940631
0.9959288059404339   0.2170217453519896   0.21456373718821004   0.38384447992245413   0.7005792004033257   0.3113682032935716   0.010828768084429095   0.4904231354313603   0.07911920456851619   0.6738017432533194   0.625134288154474   0.0018008475145853793   0.05350452170451614   0.803313400669963   0.7986590491366619   0.7024384302092032   0.7609451935596214   0.9871537212465694   0.024998616758101826   0.3967330632475946   0.04688395406698015   0.2637231923826246   0.13134235529406538   0.9833042849535315   0.050955148126546265   0.046701447030634995   0.9167786181058554   0.5994598050310774   0.35037594772322056   0.7353332437370633   0.9059498500214263   0.10903666959971711   0.2712567431547044   0.06153150048374397   0.28081556186695217   0.10723582208513174   0.21775222145018824   0.25821809981378097   0.48215651273029025   0.4047973918759286   0.4568070278905668   0.2710643785672116   0.4571578959721884   0.008064328628333972   0.40992307382358667   0.00734118618458702   0.3258155406781231   0.024760043674802446   0.35896792569704045   0.9606397391539521   0.40903692257226776   0.42530023864372507   0.008591977973819848   0.22530649541688866   0.5030870725508415   0.31626356904400793   0.7373352348191154   0.16377499493314468   0.22227151068388937   0.20902774695887621   0.5195830133689272   0.9055568951193637   0.7401149979535991   0.8042303550829476
0.06277598547836039   0.6344925165521521   0.28295710198141066   0.7961660264546137   0.6528529116547737   0.6271513303675651   0.9571415613032875   0.7714059827798112   0.29388498595773327   0.666511591213613   0.5481046387310198   0.34610574413608614   0.28529300798391344   0.4412050957967244   0.045017566180178305   0.029842175092078177   0.547957773164798   0.2774301008635797   0.822746055496289   0.8208144281332019   0.02837475979587074   0.371873205744216   0.08263105754268986   0.016584073050254364   0.9655987743175104   0.7373806891920639   0.7996739555612792   0.22041804659564074   0.31274586266273663   0.11022935882449879   0.8425323942579916   0.44901206381582953   0.018860876705003374   0.4437177676108857   0.29442775552697176   0.10290631967974342   0.7335678687210899   0.0025126718141613227   0.2494101893467935   0.07306414458766525   0.185610095556292   0.7250825709505816   0.4266641338505045   0.25224971645446326   0.15723533576042123   0.3532093652063656   0.34403307630781466   0.23566564340420892   0.19163656144291089   0.6158286760143017   0.5443591207465355   0.015247596808568183   0.8788906987801742   0.5055993171898029   0.7018267264885438   0.5662355329927387   0.8600298220751709   0.06188154957891721   0.40739897096157207   0.4633292133129952   0.12646195335408092   0.059368877764755884   0.15798878161477858   0.39026506872532996
0.9408518577977889   0.33428630681417426   0.7313246477642741   0.13801535227086667   0.7836165220373676   0.9810769416078087   0.38729157145645937   0.9023497088666578   0.5919799605944568   0.3652482655935069   0.842932450709924   0.8871021120580895   0.7130892618142826   0.859648948403704   0.14110572422138007   0.32086657906535093   0.8530594397391117   0.7977673988247868   0.733706753259808   0.8575373657523557   0.7265974863850307   0.7383985210600309   0.5757179716450294   0.4672722970270258   0.7857456285872418   0.40411221424585664   0.8443933238807554   0.3292569447561591   0.002129106549874131   0.42303527263804797   0.45710175242429596   0.42690723588950136   0.41014914595541735   0.057787007044541046   0.614169301714372   0.5398051238314118   0.6970598841411347   0.19813805864083706   0.47306357749299194   0.2189385447660608   0.844000444402023   0.40037065981605025   0.7393568242331839   0.36140117901370505   0.11740295801699228   0.6619721387560193   0.16363885258815453   0.8941288819866793   0.33165732942975046   0.2578599245101627   0.3192455287073992   0.5648719372305202   0.3295282228798763   0.8348246518721147   0.8621437762831032   0.13796470134101885   0.919379076924459   0.7770376448275736   0.24797447456873123   0.5981595775096071   0.22231919278332424   0.5788995861867366   0.7749108970757392   0.3792210327435463
0.3783187483813012   0.17852892637068637   0.03555407284255533   0.017819853729841215   0.2609157903643089   0.5165567876146671   0.8719152202544008   0.12369097174316192   0.9292584609345584   0.25869686310450435   0.5526696915470016   0.5588190345126417   0.5997302380546822   0.42387221123238966   0.6905259152638984   0.42085433317162285   0.6803511611302232   0.646834566404816   0.44255144069516716   0.8226947556620158   0.4580319683468989   0.0679349802180794   0.6676405436194279   0.4434737229184695   0.07971321996559773   0.889406053847393   0.6320864707768725   0.42565386918862824   0.8187974296012888   0.372849266232726   0.7601712505224717   0.30196289744546634   0.8895389686667303   0.11415240312822164   0.20750155897547012   0.7431438629328246   0.2898087306120482   0.690280191895832   0.5169756437115718   0.32228952976120173   0.6094575694818251   0.04344562549101598   0.07442420301640461   0.49959477409918596   0.15142560113492615   0.9755106452729366   0.4067836593969767   0.056121051180716496   0.07171238116932843   0.08610459142554354   0.7746971886201042   0.6304671819920883   0.2529149515680396   0.7132553251928175   0.014525938097632416   0.3285042845466219   0.36337598290130924   0.5991029220645959   0.8070243791221623   0.5853604216137973   0.07356725228926105   0.9088227301687639   0.2900487354105905   0.2630708918525955
0.464109682807436   0.865377104677748   0.2156245323941859   0.7634761177534095   0.31268408167250983   0.8898664594048113   0.8088408729972092   0.7073550665726931   0.2409717005031814   0.8037618679792679   0.034143684377105035   0.07688788458060482   0.9880567489351418   0.09050654278645028   0.01961774627947262   0.748383600033983   0.6246807660338325   0.4914036207218544   0.21259336715731034   0.16302317842018565   0.5511135137445715   0.5825808905530905   0.9225446317467199   0.8999522865675901   0.08700383093713548   0.7172037858753425   0.7069200993525339   0.13647616881418057   0.7743197492646257   0.8273373264705312   0.8980792263553247   0.42912110224148753   0.5333480487614443   0.02357545849126334   0.8639355419782196   0.3522332176608827   0.5452912998263024   0.9330689157048131   0.844317795698747   0.6038496176268998   0.9206105337924699   0.4416652949829587   0.6317244285414367   0.4408264392067141   0.3694970200478985   0.8590844044298682   0.7091797967947169   0.540874152639124   0.282493189110763   0.1418806185545257   0.002259697442182988   0.4043979838249434   0.5081734398461374   0.3145432920839945   0.1041804710868583   0.9752768815834559   0.9748253910846931   0.29096783359273115   0.24024492910863865   0.6230436639225732   0.4295340912583906   0.3578989178879181   0.3959271334098916   0.01919404629567343
0.5089235574659207   0.9162336229049595   0.7642027048684549   0.5783676070889593   0.1394265374180222   0.05714921847509123   0.05502290807373804   0.037493454449835296   0.8569333483072592   0.9152685999205655   0.05276321063155505   0.6330954706248919   0.34875990846112187   0.6007253078365711   0.9485827395446967   0.657818589041436   0.37393451737642874   0.30975747424383987   0.7083378104360581   0.034774925118862744   0.9444004261180382   0.9518585563559218   0.3124106770261665   0.015580878823189313   0.4354768686521175   0.03562493345096229   0.5482079721577116   0.43721327173423   0.29605033123409535   0.978475714975871   0.49318506408397356   0.3997198172843947   0.43911698292683615   0.06320711505530552   0.44042185345241847   0.7666243466595029   0.0903570744657143   0.4624818072187345   0.4918391139077217   0.10880575761806689   0.7164225570892855   0.15272433297489463   0.7835013034716636   0.07403083249920415   0.7720221309712474   0.2008657766189729   0.47109062644549715   0.05844995367601484   0.33654526231912985   0.1652408431680106   0.9228826542877856   0.6212366819417848   0.04049493108503453   0.18676512819213953   0.42969759020381204   0.22151686465739012   0.6013779481581983   0.12355801313683402   0.9892757367513936   0.45489251799788727   0.5110208736924841   0.6610762059180996   0.49743662284367185   0.3460867603798204
0.7945983166031986   0.5083518729432049   0.7139353193720082   0.2720559278806162   0.02257618563195119   0.307486096324232   0.24284469292651106   0.2136059742046014   0.6860309233128213   0.1422452531562214   0.3199620386387255   0.5923692922628165   0.6455359922277868   0.9554801249640819   0.8902644484349135   0.37085242760542647   0.044158044069588405   0.8319221118272478   0.9009887116835199   0.9159599096075391   0.5331371703771043   0.17084590590914833   0.4035520888398481   0.5698731492277188   0.7385388537739057   0.6624940329659434   0.6896167694678399   0.2978172213471026   0.7159626681419545   0.3550079366417114   0.44677207654132883   0.08421124714250117   0.029931744829133227   0.21276268348548996   0.1268100379026033   0.49184195487968463   0.38439575260134645   0.2572825585214081   0.23654558946768983   0.12098952727425816   0.34023770853175805   0.42536044669416023   0.3355568777841699   0.20502961766671898   0.8071005381546538   0.2545145407850119   0.9320047889443218   0.6351564684390002   0.06856168438074797   0.5920205078190685   0.2423880194764819   0.3373392470918976   0.3525990162387934   0.23701257117735705   0.795615942935153   0.25312799994939644   0.3226672714096602   0.02424988769186708   0.6688059050325498   0.7612860450697119   0.9382715188083137   0.766967329170459   0.4322603155648599   0.6402965177954537
0.5980338102765557   0.3416068824762988   0.09670343778069   0.4352669001287347   0.790933272121902   0.08709234169128692   0.1646986488363682   0.8001104316897345   0.7223715877411541   0.4950718338722185   0.9223106293598863   0.4627711845978369   0.3697725715023606   0.2580592626948614   0.12669468642473322   0.20964318464844042   0.047105300092700426   0.23380937500299434   0.4578887813921835   0.4483571395787286   0.10883378128438667   0.4668420458325353   0.025628465827323574   0.8080606217832749   0.5107999710078309   0.12523516335623655   0.9289250280466336   0.3727937216545402   0.7198666988859289   0.038142821664949624   0.7642263792102654   0.5726832899648057   0.997495111144775   0.5430709877927312   0.8419157498503791   0.10991210536696883   0.6277225396424143   0.28501172509786976   0.7152210634256458   0.9002689207185284   0.5806172395497139   0.051202350094875435   0.25733228203346237   0.45191178113979985   0.4717834582653272   0.5843603042623401   0.2317038162061388   0.6438511593565249   0.9609834872574963   0.45912514090610357   0.3027787881595052   0.27105743770198476   0.2411167883715673   0.4209823192411539   0.5385524089492398   0.698374147737179   0.24362167722679237   0.8779113314484228   0.6966366590988607   0.5884620423702102   0.6158991375843781   0.592899606350553   0.9814155956732149   0.6881931216516818
0.03528189803466417   0.5416972562556776   0.7240833136397525   0.23628134051188196   0.563498439769337   0.9573369519933375   0.4923794974336137   0.5924301811553571   0.6025149525118407   0.4982118110872339   0.1896007092741085   0.3213727434533723   0.3613981641402734   0.07722949184607998   0.6510483003248687   0.6229985957161932   0.11777648691348104   0.1993181603976572   0.9544116412260079   0.03453655334598304   0.501877349329103   0.6064185540471042   0.972996045552793   0.3463434316943012   0.4665954512944388   0.06472129779142662   0.24891273191304047   0.11006209118241926   0.9030970115251018   0.10738434579808914   0.7565332344794268   0.5176319100270622   0.3005820590132611   0.6091725347108552   0.5669325252053182   0.19625916657368994   0.9391838948729877   0.5319430428647752   0.9158842248804496   0.5732605708574967   0.8214074079595066   0.332624882467118   0.9614725836544417   0.5387240175115137   0.3195300586304037   0.7262063284200139   0.9884765381016487   0.1923805858172124   0.8529346073359648   0.6614850306285872   0.7395638061886082   0.08231849463479314   0.949837595810863   0.5541006848304981   0.9830305717091815   0.5646865846077309   0.6492555367976018   0.9449281501196428   0.41609804650386323   0.368427418034041   0.7100716419246141   0.4129851072548676   0.5002138216234137   0.7951668471765443
0.8886642339651075   0.08036022478774957   0.538741237968972   0.2564428296650307   0.5691341753347038   0.3541538963677357   0.5502646998673233   0.06406224384781826   0.716199567998739   0.6926688657391485   0.810700893678715   0.9817437492130251   0.7663619721878759   0.13856818090865042   0.8276703219695336   0.4170571646052942   0.11710643539027404   0.19364003078900754   0.4115722754656703   0.04862974657125323   0.40703479346565985   0.7806549235341399   0.9113584538422567   0.2534628993947089   0.5183705595005523   0.7002946987463904   0.3726172158732847   0.9970200697296783   0.9492363841658485   0.34614080237865463   0.8223525160059615   0.9329578258818599   0.23303681616710958   0.6534719366395062   0.011651622327246433   0.9512140766688348   0.46667484397923364   0.5149037557308558   0.18398130035771285   0.5341569120635407   0.3495684085889596   0.3212637249418482   0.7724090248920426   0.4855271654922874   0.9425336151232998   0.5406088014077083   0.8610505710497858   0.23206426609757852   0.4241630556227474   0.8403141026613179   0.48843335517650105   0.23504419636790025   0.4749266714568989   0.4941733002826632   0.6660808391705396   0.30208637048604026   0.24188985528978926   0.8407013636431571   0.6544292168432931   0.3508722938172054   0.7752150113105556   0.3257976079123013   0.47044791648558026   0.8167153817536648
0.425646602721596   0.004533882970453123   0.6980388915935378   0.33118821626137734   0.48311298759829624   0.46392508156274487   0.8369883205437519   0.09912395016379882   0.05894993197554882   0.623610978901427   0.3485549653672509   0.8640797537958985   0.58402326051865   0.12943767861876382   0.6824741261967113   0.5619933833098583   0.3421334052288607   0.28873631497560676   0.028044909353418187   0.21112108949265287   0.5669183939183051   0.9629387070633054   0.5575969928678379   0.3944057077389881   0.1412717911967091   0.9584048240928523   0.8595581012743001   0.06321749147761076   0.6581588035984128   0.49447974253010746   0.022569780730548154   0.964093541313812   0.5992088716228641   0.8708687636286805   0.6740148153632972   0.10001378751791339   0.015185611104214108   0.7414310850099166   0.9915406891665859   0.5380204042080551   0.6730522058753534   0.4526947700343098   0.9634957798131677   0.32689931471540223   0.10613381195704835   0.4897560629710043   0.4058987869453298   0.9324936069764141   0.9648620207603392   0.5313512388781519   0.5463406856710297   0.8692761154988033   0.3067032171619264   0.036871496348044534   0.5237709049404815   0.9051825741849915   0.7074943455390623   0.1660027327193641   0.8497560895771843   0.805168786667078   0.6923087344348482   0.4245716477094475   0.8582154004105984   0.26714838245902295
0.019256528559494775   0.9718768776751376   0.8947196205974307   0.9402490677436207   0.9131227166024465   0.4821208147041333   0.48882083365210083   0.007755460767206567   0.9482606958421071   0.9507695758259813   0.9424801479810712   0.1384793452684032   0.6415574786801808   0.9138980794779368   0.4187092430405896   0.23329677108341176   0.9340631331411186   0.7478953467585727   0.5689531534634052   0.4281279844163337   0.2417543987062703   0.3233236990491252   0.710737753052807   0.16097960195731076   0.22249787014677552   0.35144682137398753   0.8160181324553762   0.22073053421369004   0.3093751535443291   0.8693260066698542   0.3271972988032754   0.21297507344648348   0.3611144577022219   0.9185564308438728   0.38471715082220426   0.07449572817808028   0.7195569790220411   0.004658351365936092   0.9660079077816146   0.8411989570946685   0.7854938458809226   0.2567630046073634   0.39705475431820936   0.4130709726783348   0.5437394471746523   0.9334393055582382   0.6863170012654024   0.25209137072102406   0.32124157702787676   0.5819924841842506   0.8702988688100263   0.03136083650733404   0.01186642348354767   0.7126664775143965   0.5431015700067509   0.8183857630608505   0.6507519657813258   0.7941100466705235   0.1583844191845466   0.7438900348827703   0.9311949867592847   0.7894516953045875   0.19237651140293194   0.9026910777881018
0.14570114087836206   0.5326886906972241   0.7953217570847225   0.48962010510976695   0.6019616937037098   0.5992493851389858   0.10900475581932012   0.23752873438874283   0.28072011667583296   0.017256900954735217   0.23870588700929388   0.2061678978814088   0.2688536931922853   0.30459042344033876   0.6956043170025431   0.38778213482055823   0.6181017274109596   0.5104803767698152   0.5372198978179965   0.643892099937788   0.6869067406516749   0.7210286814652277   0.3448433864150645   0.7412010221496862   0.5412055997733128   0.1883399907680036   0.549521629330342   0.25158091703991925   0.9392439060696031   0.5890906056290177   0.44051687351102187   0.01405218265117643   0.6585237893937701   0.5718337046742825   0.20181098650172796   0.8078842847697676   0.3896700962014848   0.26724328123394375   0.5062066694991849   0.4201021499492094   0.7715683687905253   0.7567629044641285   0.9689867716811884   0.7762100500114215   0.08466162813885034   0.035734222998900896   0.6241433852661239   0.03500902786173527   0.5434560283655375   0.8473942322308973   0.07462175593578194   0.783428110821816   0.6042121222959344   0.2583036266018796   0.63410488242476   0.7693759281706396   0.9456883329021643   0.6864699219275971   0.43229389592303213   0.9614916434008719   0.5560182367006794   0.41922664069365345   0.9260872264238472   0.5413894934516625
0.7844498679101541   0.6624637362295248   0.9571004547426588   0.765179443440241   0.6997882397713038   0.626729513230624   0.3329570694765349   0.7301704155785058   0.15633221140576636   0.7793352809997267   0.258335313540753   0.9467423047566897   0.552120089109832   0.521031654397847   0.6242304311159929   0.17736637658605023   0.6064317562076678   0.8345617324702499   0.19193653519296075   0.21587473318517827   0.05041351950698833   0.41533509177659644   0.2658493087691135   0.6744852397335157   0.26596365159683416   0.7528713555470715   0.3087488540264547   0.9093057962932747   0.5661754118255303   0.1261418423164476   0.9757917845499198   0.17913538071476887   0.40984320041976396   0.34680656131672094   0.7174564710091668   0.23239307595807907   0.857723111309932   0.8257749069188739   0.09322603989317389   0.05502669937202885   0.25129135510226425   0.991213174448624   0.9012895047002132   0.8391519661868506   0.20087783559527592   0.5758780826720276   0.6354401959310997   0.16466672645333483   0.9349141839984417   0.823006727124956   0.32669134190464494   0.2553609301600602   0.3687387721729114   0.6968648848085084   0.3508995573547252   0.0762255494452913   0.9588955717531474   0.3500583234917875   0.6334430863455585   0.8438324734872122   0.10117246044321546   0.5242834165729136   0.5402170464523846   0.7888057741151834
0.8498811053409512   0.5330702421242896   0.6389275417521714   0.9496538079283328   0.6490032697456753   0.957192159452262   0.003487345821071736   0.784987081474998   0.7140890857472336   0.13418543232730593   0.6767960039164268   0.5296261513149378   0.34535031357432217   0.4373205475187975   0.3258964465617016   0.4534006018696465   0.38645474182117473   0.08726222402701003   0.6924533602161431   0.6095681283824342   0.28528228137795925   0.5629788074540965   0.15223631376375865   0.820762354267251   0.43540117603700806   0.029908565329806926   0.5133087720115873   0.8711085463389181   0.7863979062913328   0.07271640587754498   0.5098214261905155   0.08612146486392017   0.07230882054409915   0.9385309735502391   0.8330254222740887   0.5564953135489824   0.726958506969777   0.5012104260314415   0.5071289757123871   0.10309471167933587   0.3405037651486023   0.4139482020044315   0.814675615496244   0.4935265832969016   0.05522148377064303   0.850969394550335   0.6624393017324853   0.6727642290296507   0.619820307733635   0.8210608292205281   0.1491305297208981   0.8016556826907325   0.8334224014423023   0.7483444233429831   0.6393091035303826   0.7155342178268124   0.7611135808982031   0.8098134497927441   0.8062836812562938   0.15903890427783   0.03415507392842611   0.30860302376130255   0.29915470554390666   0.05594419259849411
0.6936513087798238   0.894654821756871   0.48447909004766265   0.5624176093015926   0.6384298250091808   0.043685427206536   0.8220397883151773   0.8896533802719419   0.018609517275545787   0.2226245979860079   0.6729092585942792   0.0879976975812093   0.18518711583324352   0.47428017464302474   0.03360015506389663   0.3724634797543969   0.4240735349350404   0.6644667248502807   0.2273164738076028   0.21342457547656693   0.3899184610066143   0.35586370108897813   0.9281617682636961   0.1574803828780728   0.6962671522267905   0.4612088793321071   0.44368267821603347   0.5950627735764803   0.05783732721760971   0.41752345212557107   0.6216428899008561   0.7054093933045384   0.03922780994206392   0.19489885413956318   0.948733631306577   0.6174116957233291   0.8540406941088204   0.7206186794965385   0.9151334762426804   0.24494821596893224   0.42996715917378   0.05615195464625775   0.6878170024350776   0.03152364049236529   0.040048698167165685   0.7002882535572796   0.7596552341713814   0.8740432576142925   0.3437815459403752   0.23907937422517256   0.3159725559553479   0.27898048403781217   0.2859442187227655   0.8215559220996015   0.6943296660544918   0.5735710907332737   0.24671640878070156   0.6266570679600383   0.7455960347479148   0.9561593950099445   0.39267571467188117   0.9060383884634999   0.8304625585052344   0.7112111790410124
0.9627085554981012   0.8498864338172422   0.1426455560701569   0.679687538548647   0.9226598573309355   0.14959818025996252   0.38299032189877547   0.8056442809343546   0.5788783113905603   0.91051880603479   0.06701776594342754   0.5266637968965424   0.2929340926677948   0.08896288393518845   0.3726880998889358   0.9530927061632687   0.046217683887093235   0.46230581597515014   0.627092065141021   0.9969333111533242   0.6535419692152121   0.5562674275116503   0.7966295066357866   0.2857221321123118   0.6908334137171109   0.7063809936944081   0.6539839505656297   0.6060345935636647   0.7681735563861755   0.5567828134344456   0.2709936286668543   0.8003903126293102   0.18929524499561515   0.6462640073996556   0.20397586272342672   0.2737265157327678   0.8963611523278203   0.5573011234644671   0.8312877628344909   0.3206338095694991   0.8501434684407271   0.09499530748931703   0.2041956976934699   0.32370049841617493   0.19660149922551504   0.5387278799776668   0.40756619105768327   0.03797836630386317   0.5057680855084041   0.8323468862832587   0.7535822404920536   0.4319437727401984   0.7375945291222287   0.2755640728488132   0.4825886118251993   0.6315534601108883   0.5482992841266136   0.6293000654491576   0.2786127491017726   0.3578269443781205   0.6519381317987932   0.07199894198469044   0.4473249862672816   0.03719313480862141
0.8017946633580662   0.9770036344953734   0.24312928857381175   0.7134926363924464   0.6051931641325511   0.4382757545177066   0.8355630975161285   0.6755142700885832   0.09942507862414698   0.6059288682344479   0.08198085702407491   0.24357049734838485   0.3618305495019183   0.3303647953856347   0.5993922451988756   0.6120170372374966   0.8135312653753047   0.7010647299364771   0.32077949609710305   0.2541900928593761   0.16159313357651148   0.6290657879517867   0.8734545098298214   0.2169969580507547   0.35979847021844535   0.6520621534564133   0.6303252212560096   0.5035043216583083   0.7546053060858943   0.21378639893870666   0.7947621237398812   0.8279900515697249   0.6551802274617473   0.6078575307042587   0.7127812667158063   0.5844195542213401   0.29334967795982897   0.2774927353186241   0.1133890215169307   0.9724025169838435   0.47981841258452423   0.576428005382147   0.7926095254198277   0.7182124241244674   0.3182252790080128   0.9473622174303603   0.9191550155900062   0.5012154660737127   0.9584268087895674   0.2953000639739471   0.2888297943339965   0.9977111444154044   0.20382150270367316   0.08151366503524045   0.49406767059411527   0.1697210928456795   0.5486412752419259   0.47365613433098164   0.7812864038783089   0.5853015386243394   0.25529159728209694   0.19616339901235755   0.6678973823613783   0.6128990216404958
0.7754731846975726   0.6197353936302106   0.8752878569415506   0.8946865975160284   0.45724790568955986   0.6723731761998502   0.9561328413515444   0.3934711314423157   0.4988210968999925   0.37707311222590306   0.667303047017548   0.39575998702691123   0.2949995941963193   0.2955594471906626   0.17323537642343265   0.22603889418123174   0.7463583189543934   0.821903312859681   0.39194897254512373   0.6407373555568924   0.49106672167229654   0.6257399138473234   0.7240515901837454   0.027838333916396528   0.7155935369747238   0.006004520217112896   0.8487637332421949   0.1331517364003681   0.25834563128516397   0.3336313440172627   0.8926308918906504   0.7396806049580524   0.7595245343851715   0.9565582317913596   0.2253278448731025   0.34392061793114115   0.46452494018885215   0.6609987846006969   0.05209246844966983   0.11788172374990938   0.7181666212344587   0.839095471741016   0.6601434959045461   0.477144368193017   0.22709989956216223   0.21335555789369257   0.9360919057208007   0.44930603427662047   0.5115063625874384   0.20735103767657967   0.0873281724786058   0.3161542978762524   0.2531607313022744   0.8737196936593169   0.19469728058795538   0.5764736929181999   0.4936361969171029   0.9171614618679573   0.9693694357148529   0.23255307498705885   0.029111256728250743   0.25616267726726033   0.917276967265183   0.11467135123714947
0.310944635493792   0.4170672055262444   0.2571334713606369   0.6375269830441325   0.08384473593162976   0.2037116476325518   0.32104156563983627   0.188220948767512   0.5723383733441914   0.9963606099559721   0.2337133931612305   0.8720666508912597   0.31917764204191695   0.12264091629665519   0.03901611257327511   0.2955929579730596   0.8255414451248141   0.20547945442869786   0.06964667685842221   0.06303988298600077   0.7964301883965633   0.9493167771614375   0.15236970959323917   0.9483685317488513   0.4854855529027713   0.5322495716351932   0.8952362382326022   0.3108415487047188   0.40164081697114157   0.3285379240026413   0.5741946725927659   0.12262059993720684   0.8293024436269502   0.3321773140466692   0.34048127943153544   0.2505539490459472   0.5101248015850331   0.209536397750014   0.30146516685826036   0.9549609910728876   0.6845833564602192   0.0040569433213161615   0.23181848999983815   0.8919211080868868   0.8881531680636559   0.05474016615987866   0.07944878040659897   0.9435525763380355   0.40266761516088456   0.5224905945246855   0.18421254217399674   0.6327110276333167   0.0010267981897429937   0.19395267052204418   0.6100178695812308   0.5100904276961098   0.1717243545627928   0.861775356475375   0.26953659014969533   0.2595364786501626   0.6615995529777596   0.652238958725361   0.968071423291435   0.30457548757727504
0.9770161965175405   0.6481820154040449   0.7362529332915968   0.41265437949038825   0.08886302845388461   0.5934418492441661   0.6568041528849978   0.4691018031523528   0.686195413293   0.07095125471948062   0.47259161071100114   0.8363907755190361   0.6851686151032571   0.8769985841974365   0.8625737411297704   0.3263003478229263   0.5134442605404642   0.015223227722061453   0.593037150980075   0.06676386917276364   0.8518447075627046   0.3629842689967005   0.62496572768864   0.7621883815954886   0.8748285110451641   0.7148022535926557   0.8887127943970432   0.3495340021051003   0.7859654825912795   0.12136040434848952   0.23190864151204532   0.8804321989527476   0.0997700692982795   0.0504091496290089   0.7593170308010442   0.04404142343371147   0.4146014541950224   0.17341056543157246   0.8967432896712738   0.7177410756107853   0.9011571936545582   0.15818733770951102   0.30370613869119883   0.6509772064380216   0.04931248609185355   0.7952030687128105   0.6787404110025588   0.888788824842533   0.1744839750466894   0.08040081512015484   0.7900276166055156   0.5392548227374326   0.3885184924554098   0.9590404107716654   0.5581189750934702   0.6588226237846851   0.28874842315713034   0.9086312611426565   0.798801944292426   0.6147812003509736   0.8741469689621079   0.735220695711084   0.9020586546211522   0.8970401247401883
0.9729897753075497   0.577033358001573   0.5983525159299534   0.24606291830216684   0.9236772892156961   0.7818302892887624   0.9196121049273946   0.35727409345963385   0.7491933141690068   0.7014294741686076   0.12958448832187908   0.8180192707222012   0.360674821713597   0.7423890633969422   0.5714655132284089   0.15919664693751606   0.07192639855646665   0.8337578022542859   0.7726635689359828   0.5444154465865425   0.19777942959435876   0.09853710654320186   0.8706049143148306   0.647375321846354   0.22478965428680905   0.5215037485416288   0.2722523983848772   0.40131240354418724   0.3011123650711129   0.7396734592528664   0.35264029345748255   0.044038310084553396   0.5519190509021061   0.03824398508425885   0.22305580513560347   0.22601903936235224   0.19124422918850917   0.2958549216873166   0.6515902919071946   0.06682239242483616   0.1193178306320425   0.4620971194330308   0.8789267229712118   0.5224069458382937   0.9215384010376837   0.36356001288982887   0.008321808656381203   0.8750316239919397   0.6967487467508746   0.8420562643482   0.736069410271504   0.47371922044775244   0.3956363816797618   0.10238280509533355   0.3834291168140215   0.42968091036319905   0.8437173307776556   0.0641388200110747   0.16037331167841798   0.2036618710008468   0.6524731015891465   0.7682838983237581   0.5087830197712234   0.13683947857601064
0.533155270957104   0.3061867788907274   0.6298562968000115   0.6144325327377169   0.6116168699194202   0.9426267660008985   0.6215344881436303   0.7394009087457774   0.9148681231685456   0.10057050165269847   0.8854650778721264   0.26568168829802485   0.5192317414887838   0.998187696557365   0.5020359610581049   0.8360007779348259   0.6755144107111282   0.9340488765462902   0.34166264937968693   0.6323389069339791   0.023041309121981695   0.1657649782225321   0.8328796296084635   0.4954994283579684   0.4898860381648777   0.8595781993318048   0.20302333280845197   0.8810668956202514   0.8782691682454574   0.9169514333309063   0.5814888446648216   0.14166598687447415   0.9634010450769118   0.8163809316782078   0.6960237667926953   0.8759842985764492   0.44416930358812806   0.8181932351208429   0.19398780573459035   0.03998352064162342   0.7686548928769998   0.8841443585745526   0.8523251563549035   0.4076446137076444   0.7456135837550182   0.7183793803520205   0.019445526746439887   0.912145185349676   0.2557275455901405   0.8588011810202159   0.8164221939379879   0.031078289729424544   0.377458377344683   0.9418497476893095   0.2349333492731663   0.8894123028549504   0.41405733226777114   0.1254688160111017   0.538909582480471   0.013428004278501125   0.9698880286796431   0.3072755808902588   0.3449217767458807   0.9734444836368777
0.2012331358026432   0.4231312223157061   0.4925966203909773   0.5657998699292334   0.45561955204762505   0.7047518419636856   0.4731510936445374   0.6536546845795573   0.19989200645748456   0.8459506609434697   0.6567288997065495   0.6225763948501328   0.8224336291128016   0.9041009132541602   0.4217955504333832   0.7331640919951824   0.4083762968450304   0.7786320972430585   0.8828859679529121   0.7197360877166813   0.43848826816538733   0.4713565163527997   0.5379641912070314   0.7462916040798035   0.2372551323627441   0.04822529403709356   0.045367570816054165   0.18049173415057024   0.781635580315119   0.343473452073408   0.5722164771715168   0.526837049571013   0.5817435738576345   0.4975227911299383   0.9154875774649673   0.9042606547208801   0.7593099447448329   0.593421877875778   0.49369202703158416   0.17109656272569773   0.3509336478998026   0.8147897806327197   0.610806059078672   0.4513604750090165   0.9124453797344152   0.34343326427991994   0.07284186787164058   0.7050688709292129   0.6751902473716711   0.29520797024282636   0.027474297055586423   0.5245771367786427   0.8935546670565521   0.9517345181694183   0.45525781988406966   0.9977400872076297   0.31181109319891753   0.45421172703948004   0.5397702424191023   0.09347943248674961   0.5525011484540846   0.8607898491637019   0.046078215387518176   0.9223828697610519
0.20156750055428205   0.04600006853098234   0.43527215630884614   0.4710223947520354   0.2891221208198668   0.7025668042510624   0.3624302884372056   0.7659535238228226   0.6139318734481957   0.407358834008236   0.33495599138161913   0.24137638704417985   0.7203772063916436   0.4556243158388177   0.8796981714975495   0.2436362998365501   0.40856611319272607   0.0014125887993376033   0.3399279290784472   0.1501568673498005   0.8560649647386415   0.14062273963563565   0.293849713690929   0.2277739975887486   0.6544974641843594   0.0946226711046533   0.8585775573820829   0.7567516028367132   0.3653753433644926   0.3920558668535909   0.49614726894487726   0.9907980790138907   0.751443469916297   0.9846970328453549   0.16119127756325813   0.7494216919697109   0.031066263524653352   0.5290727170065372   0.2814931060657086   0.5057853921331608   0.6225001503319273   0.5276601282071997   0.9415651769872614   0.35562852478336027   0.7664351855932858   0.38703738857156395   0.6477154632963324   0.12785452719461163   0.11193772140892644   0.29241471746691067   0.7891379059142496   0.3711029243578984   0.7465623780444338   0.9003588506133198   0.2929906369693723   0.3803048453440077   0.9951189081281369   0.9156618177679648   0.13179935940611417   0.6308831533742969   0.9640526446034835   0.38658910076142766   0.8503062533404055   0.1250977612411361
0.3415524942715562   0.8589289725542281   0.9087410763531442   0.7694692364577759   0.5751173086782704   0.4718915839826641   0.2610256130568117   0.6416147092631642   0.4631795872693439   0.17947686651575345   0.4718877071425621   0.27051178490526584   0.7166172092249101   0.2791180159024337   0.17889707017318981   0.8902069395612582   0.7214983010967732   0.36345619813446883   0.04709771076707565   0.2593237861869613   0.7574456564932897   0.9768670973730411   0.1967914574266701   0.1342260249458252   0.41589316222173345   0.11793812481881305   0.288050381073526   0.3647567884880493   0.8407758535434631   0.6460465408361489   0.0270247680167143   0.723142079224885   0.3775962662741192   0.4665696743203955   0.5551370608741522   0.4526302943196192   0.6609790570492091   0.18745165841796177   0.37623999070096237   0.5624233547583611   0.939480755952436   0.8239954602834929   0.32914227993388673   0.3030995685713998   0.18203509945914623   0.8471283629104518   0.1323508225072166   0.1688735436255746   0.7661419372374128   0.7291902380916387   0.8443004414336907   0.8041167551375252   0.9253660836939497   0.08314369725548984   0.8172756734169764   0.08097467591264021   0.5477698174198304   0.6165740229350943   0.2621386125428241   0.628344381593021   0.8867907603706213   0.4291223645171326   0.8858986218418617   0.06592102683465989
0.9473100044181854   0.6051269042336397   0.5567563419079751   0.7628214582632601   0.7652749049590392   0.7579985413231879   0.42440551940075844   0.5939479146376855   0.9991329677216264   0.02880830323154908   0.5801050779670678   0.7898311595001603   0.07376688402767674   0.9456646059760593   0.7628294045500915   0.70885648358752   0.5259970666078463   0.32909058304096483   0.5006907920072673   0.08051210199449903   0.639206306237225   0.8999682185238322   0.6147921701654055   0.014591075159839144   0.6918963018190396   0.29484131429019256   0.058035828257430526   0.25176961689657906   0.9266213968600004   0.5368427729670048   0.6336303088566722   0.6578217022588936   0.927488429138374   0.5080344697354556   0.0535252308896043   0.8679905427587333   0.8537215451106973   0.5623698637593965   0.29069582633951285   0.15913405917121332   0.32772447850285097   0.23327928071843154   0.7900050343322454   0.07862195717671429   0.6885181722656261   0.33331106219459933   0.17521286416683993   0.06403088201687515   0.9966218704465865   0.038469747904406736   0.1171770359094094   0.8122612651202961   0.07000047358658607   0.501626974937402   0.48354672705273727   0.15443956286140256   0.14251204444821206   0.9935925052019463   0.430021496163133   0.2864490201026692   0.28879049933751477   0.43122264144254996   0.13932566982362016   0.1273149609314559
0.9610660208346639   0.1979433607241184   0.34932063549137465   0.048693003754741615   0.2725478485690378   0.8646322985295191   0.17410777132453475   0.9846621217378665   0.27592597812245134   0.8261625506251123   0.05693073541512536   0.17240085661757037   0.20592550453586528   0.32453557568771035   0.5733840083623881   0.017961293756167816   0.06341346008765321   0.330943070485764   0.14336251219925508   0.7315122736534986   0.7746229607501384   0.899720429043214   0.004036842375634923   0.6041973127220427   0.8135569399154746   0.7017770683190956   0.6547162068842602   0.5555043089673011   0.5410090913464368   0.8371447697895765   0.4806084355597255   0.5708421872294346   0.2650831132239855   0.010982219164464216   0.42367770014460016   0.39844133061186426   0.0591576086881202   0.6864466434767539   0.850293691782212   0.3804800368556964   0.995744148600467   0.3555035729909899   0.706931179582957   0.6489677632021978   0.22112118785032858   0.45578314394777586   0.7028943372073221   0.04477045048015514   0.407564247934854   0.7540060756286803   0.04817813032306181   0.4892661415128541   0.8665551565884172   0.9168613058391036   0.5675696947633363   0.9184239542834195   0.6014720433644317   0.9058790866746395   0.14389199461873617   0.5199826236715552   0.5423144346763116   0.21943244319788557   0.2935983028365241   0.13950258681585878
0.5465702860758446   0.8639288702068957   0.5866671232535671   0.49053482361366096   0.32544909822551593   0.4081457262591198   0.883772786046245   0.4457643731335058   0.9178848502906619   0.6541396506304396   0.8355946557231833   0.9564982316206517   0.051329693702244765   0.7372783447913359   0.2680249609598469   0.038074277337232294   0.44985765033781305   0.8313992581166965   0.12413296634111075   0.5180916536656771   0.9075432156615015   0.6119668149188109   0.8305346635045867   0.3785890668498183   0.36097292958565697   0.7480379447119152   0.24386754025101956   0.8880542432361573   0.035523831360141034   0.33989221845279544   0.3600947542047745   0.44228987010265153   0.11763898106947908   0.6857525678223558   0.5245000984815913   0.4857916384819998   0.06630928736723432   0.9484742230310199   0.2564751375217444   0.4477173611447675   0.6164516370294213   0.11707496491432347   0.13234217118063363   0.9296257074790905   0.7089084213679198   0.5051081499955126   0.30180750767604697   0.5510366406292722   0.3479354917822628   0.7570702052835974   0.05793996742502742   0.6629823973931148   0.31241166042212176   0.41717798683080193   0.697845213220253   0.22069252729046324   0.19477267935264267   0.731425419008446   0.1733451147386616   0.7349008888084635   0.12846339198540838   0.7829511959774261   0.9168699772169172   0.2871835276636959
0.512011754955987   0.6658762310631027   0.7845278060362836   0.3575578201846055   0.8031033335880673   0.1607680810675901   0.4827202983602366   0.8065211795553334   0.45516784180580455   0.40369787578399274   0.4247803309352092   0.14353878216221866   0.14275618138368276   0.9865198889531908   0.7269351177149563   0.9228462548717554   0.9479835020310401   0.2550944699447447   0.5535900029762947   0.18794536606329199   0.8195201100456317   0.4721432739673186   0.6367200257593775   0.900761838399596   0.30750835508964464   0.8062670429042159   0.8521922197230939   0.5432040182149905   0.5044050215015773   0.6454989618366258   0.3694719213628573   0.7366828386596571   0.04923717969577279   0.24180108605263304   0.944691590427648   0.5931440564974384   0.9064809983120901   0.25528119709944225   0.21775647271269175   0.670297801625683   0.95849749628105   0.00018672715469749942   0.664166469736397   0.48235243556239105   0.13897738623541822   0.5280434531873789   0.02744644397701957   0.581590597162795   0.8314690311457736   0.7217764102831631   0.1752542242539257   0.03838657894780448   0.3270640096441963   0.07627744844653726   0.8057823028910684   0.3017037402881474   0.2778268299484235   0.8344763623939042   0.8610907124634204   0.708559683790709   0.37134583163633345   0.579195165294462   0.6433342397507287   0.038261882165025934
0.41284833535528354   0.5790084381397645   0.9791677700143316   0.5559094466026349   0.2738709491198653   0.050964984952385564   0.9517213260373121   0.9743188494398399   0.44240191797409173   0.3291885746692225   0.7764671017833863   0.9359322704920354   0.11533790832989545   0.25291112622268525   0.970684798892318   0.634228530203888   0.837511078381472   0.41843476382878103   0.10959408642889752   0.9256688464131791   0.4661652467451385   0.8392395985343191   0.4662598466781689   0.8874069642481531   0.053316911389854976   0.2602311603945546   0.48709207666383725   0.33149751764551827   0.7794459622699896   0.209266175442169   0.5353707506265253   0.35717866820567834   0.33704404429589796   0.8800776007729465   0.7589036488431389   0.4212463977136429   0.22170613596600253   0.6271664745502612   0.788218849950821   0.7870178675097549   0.38419505758453054   0.20873171072148014   0.6786247635219235   0.8613490210965757   0.9180298108393921   0.3694921121871611   0.2123649168437546   0.9739420568484226   0.8647128994495371   0.10926095179260654   0.7252728401799173   0.6424445392029043   0.08526693717954742   0.8999947763504376   0.1899020895533921   0.28526587099722595   0.7482228928836494   0.01991717557749109   0.4309984407102532   0.8640194732835831   0.526516756917647   0.39275070102722986   0.6427795907594323   0.07700160577382817
0.14232169933311636   0.18401899030574975   0.9641548272375087   0.2156525846772524   0.2242918884937243   0.8145268781185886   0.7517899103937541   0.24171052782882985   0.3595789890441872   0.7052659263259821   0.026517070213836764   0.5992659886259255   0.2743120518646398   0.8052711499755446   0.8366149806604447   0.31400011762869956   0.5260891589809903   0.7853539743980534   0.4056165399501915   0.44998064434511653   0.9995724020633434   0.39260327337082357   0.7628369491907593   0.3729790385712884   0.8572507027302271   0.20858428306507382   0.7986821219532505   0.15732645389403596   0.6329588142365027   0.39405740494648517   0.046892211559496445   0.9156159260652061   0.2733798251923155   0.688791478620503   0.020375141345659684   0.3163499374392806   0.9990677733276757   0.8835203286449586   0.18376016068521503   0.002349819810581023   0.47297861434668537   0.09816635424690505   0.7781436207350235   0.5523691754654645   0.47340621228334195   0.7055630808760814   0.015306671544264286   0.17939013689417613   0.6161555095531149   0.4969787978110076   0.21662454959101374   0.022063683000140166   0.9831966953166121   0.10292139286452247   0.1697323380315173   0.10644775693493405   0.7098168701242967   0.4141299142440194   0.1493571966858576   0.7900978194956535   0.710749096796621   0.5306095855990609   0.9655970360006426   0.7877479996850725
0.2377704824499356   0.43244323135215584   0.18745341526561904   0.23537882421960796   0.7643642701665936   0.7268801504760743   0.17214674372135474   0.05598868732543182   0.1482087606134787   0.2299013526650667   0.955522194130341   0.033925004325291656   0.16501206529686652   0.12697995980054422   0.7857898560988237   0.9274772473903576   0.45519519517256984   0.7128500455565249   0.6364326594129661   0.13737942789470417   0.7444460983759489   0.18224045995746396   0.6708356234123235   0.3496314282096317   0.5066756159260133   0.7497972286053082   0.4833822081467045   0.1142526039900238   0.7423113457594197   0.022917078129233805   0.3112354644253498   0.058263916664591964   0.5941025851459409   0.7930157254641671   0.35571327029500877   0.024338912339300304   0.4290905198490744   0.6660357656636229   0.5699234141961851   0.09686166494894269   0.9738953246765045   0.953185720107098   0.9334907547832189   0.9594822370542385   0.22944922630055567   0.770945260149634   0.26265513137089536   0.6098508088446069   0.7227736103745424   0.021148031544325922   0.7792729232241908   0.495598204854583   0.9804622646151228   0.9982309534150922   0.46803745879884107   0.43733428818999104   0.38635967946918176   0.205215227950925   0.11232418850383234   0.41299537585069074   0.9572691596201074   0.5391794622873022   0.5424007743076473   0.3161337109017481
0.9833738349436029   0.5859937421802041   0.6089100195244284   0.3566514738475095   0.7539246086430471   0.81504848203057   0.346254888153533   0.7468006650029028   0.03115099826850479   0.7939004504862441   0.5669819649293422   0.2512024601483197   0.05068873365338207   0.795669497071152   0.09894450613050107   0.8138681719583287   0.6643290541842003   0.590454269120227   0.9866203176266687   0.40087279610763793   0.7070598945640929   0.05127480683292484   0.4442195433190214   0.08473908520588988   0.72368605962049   0.46528106465272073   0.835309523794593   0.7280876113583804   0.9697614509774429   0.6502325826221507   0.48905463564106   0.9812869463554776   0.9386104527089382   0.8563321321359066   0.9220726707117178   0.7300844862071579   0.8879217190555561   0.06066263506475463   0.8231281645812167   0.9162163142488292   0.22359266487135576   0.47020836594452764   0.836507846954548   0.5153435181411913   0.5165327703072629   0.4189335591116028   0.3922883036355266   0.43060443293530143   0.7928467106867728   0.9536524944588821   0.5569787798409336   0.7025168215769211   0.8230852597093299   0.30341991183673134   0.06792414419987355   0.7212298752214434   0.8844748070003917   0.44708777970082475   0.14585147348815572   0.9911453890142855   0.9965530879448358   0.38642514463607014   0.32272330890693895   0.07492907476545628
0.77296042307348   0.9162167786915425   0.4862154619523909   0.559585556624265   0.2564276527662171   0.49728321957993965   0.0939271583168643   0.12898112368896358   0.4635809420794443   0.5436307251210576   0.5369483784759307   0.4264643021120425   0.6404956823701144   0.2402108132843262   0.46902423427605716   0.7052344268905991   0.7560208753697226   0.7931230335835014   0.32317276078790147   0.7140890378763136   0.759467787424887   0.40669788894743136   0.0004494518809625284   0.6391599631108573   0.986507364351407   0.49048111025588886   0.5142339899285716   0.0795744064865923   0.7300797115851899   0.9931978906759492   0.42030683161170734   0.9505932827976288   0.2664987695057456   0.4495671655548917   0.8833584531357767   0.5241289806855862   0.6260030871356311   0.20935635227056548   0.41433421885971944   0.8188945537949871   0.8699822117659085   0.41623331868706404   0.091161458071818   0.10480551591867356   0.11051442434102157   0.009535429739632676   0.09071200619085547   0.4656455528078163   0.12400705998961462   0.5190543194837438   0.5764780162622838   0.38607114632122397   0.3939273484044248   0.5258564288077946   0.1561711846505765   0.43547786352359524   0.1274285788986792   0.07628926325290288   0.27281273151479984   0.9113488828380091   0.5014254917630481   0.8669329109823374   0.8584785126550805   0.0924543290430219
0.6314432799971396   0.4506995922952734   0.7673170545832624   0.9876488131243484   0.520928855656118   0.4411641625556407   0.676605048392407   0.5220032603165321   0.3969217956665034   0.9221098430718969   0.10012703213012313   0.13593211399530808   0.0029944472620786096   0.3962534142641024   0.9439558474795466   0.7004542504717128   0.8755658683633994   0.3199641510111995   0.6711431159647467   0.7891053676337039   0.3741403766003514   0.4530312400288621   0.8126646033096664   0.6966510385906819   0.7426970966032118   0.002331647733588716   0.045347548726403945   0.7090022254663336   0.2217682409470938   0.561167485177948   0.36874250033399697   0.18699896514980155   0.8248464452805905   0.6390576421060511   0.2686154682038739   0.05106685115449345   0.8218519980185118   0.24280422784194874   0.32465962072432725   0.3506126006827806   0.9462861296551124   0.9228400768307492   0.6535165047595805   0.5615072330490768   0.5721457530547611   0.4698088368018872   0.8408519014499141   0.8648561944583949   0.8294486564515493   0.46747718906829844   0.7955043527235102   0.15585396899206125   0.6076804155044555   0.9063097038903505   0.4267618523895132   0.9688550038422598   0.782833970223865   0.26725206178429933   0.1581463841856393   0.9177881526877663   0.9609819722053532   0.024447833942350585   0.8334867634613121   0.5671755520049857
0.014695842550240779   0.10160775711160133   0.1799702587017316   0.005668318955908882   0.4425500894954797   0.6317989203097142   0.3391183572518175   0.14081212449751404   0.6131014330439304   0.16432173124141575   0.5436140045283073   0.9849581555054527   0.005421017539474966   0.2580120273510653   0.11685215213879414   0.016103151663193056   0.22258704731560994   0.9907599655667659   0.9587057679531549   0.09831499897542678   0.2616050751102567   0.9663121316244154   0.12521900449184276   0.5311394469704411   0.24690923256001596   0.864704374512814   0.9452487457901112   0.5254711280145322   0.8043591430645363   0.23290545420309988   0.6061303885382937   0.3846590035170182   0.19125771002060582   0.06858372296168415   0.06251638400998635   0.3997008480115654   0.18583669248113086   0.8105716956106188   0.9456642318711922   0.3835976963483724   0.9632496451655209   0.8198117300438529   0.9869584639180373   0.2852826973729456   0.7016445700552641   0.8534995984194375   0.8617394594261946   0.7541432504025045   0.4547353374952482   0.9887952239066234   0.9164907136360835   0.22867212238797224   0.6503761944307119   0.7558897697035235   0.31036032509778977   0.844013118870954   0.45911848441010616   0.6873060467418394   0.24784394108780342   0.44431227085938857   0.2732817919289753   0.8767343511312206   0.3021797092166112   0.060714574511016195
0.31003214676345436   0.05692262108736766   0.3152212452985738   0.7754318771380706   0.6083875767081902   0.2034230226679302   0.4534817858723792   0.021288626735566123   0.153652239212942   0.2146277987613068   0.5369910722362958   0.7926165043475939   0.5032760447822301   0.45873802905778327   0.226630747138506   0.9486033854766399   0.04415756037212389   0.7714319823159439   0.9787868060507026   0.5042911146172513   0.7708757684431486   0.8946976311847235   0.6766070968340914   0.4435765401062351   0.4608436216796942   0.8377750100973558   0.3613858515355176   0.6681446629681645   0.852456044971504   0.6343519874294256   0.9079040656631384   0.6468560362325984   0.6988038057585619   0.4197241886681187   0.3709129934268426   0.8542395318850045   0.19552776097633193   0.9609861596103354   0.14428224628833658   0.9056361464083647   0.15137020060420803   0.18955417729439153   0.165495440237634   0.4013450317911133   0.38049443216105944   0.2948565461096681   0.48888834340354254   0.9577684916848782   0.9196508104813652   0.4570815360123124   0.12750249186802495   0.2896238287167137   0.06719476550986127   0.8227295485828868   0.21959842620488657   0.6427677924841153   0.36839095975129926   0.4030053599147681   0.848685432778044   0.7885282605991109   0.17286319877496736   0.44201920030443265   0.7044031864897073   0.8828921141907462
0.021492998170759312   0.25246502301004115   0.5389077462520734   0.4815470823996329   0.6409985660096998   0.957608476900373   0.050019402848530826   0.5237785907147546   0.7213477555283346   0.5005269408880606   0.9225169109805059   0.23415476199804097   0.6541529900184734   0.6777973923051738   0.7029184847756194   0.5913869695139257   0.28576203026717406   0.2747920323904056   0.8542330519975754   0.8028587089148148   0.11289883149220671   0.832772832085973   0.14982986550786798   0.9199665947240686   0.0914058333214474   0.5803078090759318   0.6109221192557946   0.43841951232443566   0.4504072673117475   0.6226993321755588   0.5609027164072637   0.914640921609681   0.7290595117834129   0.12217239128749824   0.6383858054267579   0.68048615961164   0.07490652176493956   0.44437499898232447   0.9354673206511386   0.08909919009771441   0.7891444914977656   0.16958296659191885   0.08123426865356324   0.28624048118289963   0.6762456600055587   0.3368101345059459   0.9314044031456953   0.3662738864588311   0.5848398266841114   0.756502325430014   0.32048228388990063   0.9278543741343954   0.13443255937236387   0.1338029932544552   0.7595795674826369   0.013213452524714387   0.40537304758895093   0.011630601966956963   0.12119376205587898   0.33272729291307435   0.33046652582401137   0.5672556029846325   0.18572644140474037   0.24362810281535993
0.5413220343262459   0.3976726363927136   0.10449217275117713   0.9573876216324603   0.8650763743206871   0.06086250188676774   0.1730877696054819   0.5911137351736293   0.2802365476365757   0.3043601764567537   0.8526054857155813   0.6632593610392339   0.14580398826421181   0.17055718320229848   0.09302591823294434   0.6500459085145195   0.7404309406752608   0.15892658123534154   0.9718321561770654   0.31731861560144514   0.4099644148512495   0.591670978250709   0.786105714772325   0.0736905127860852   0.8686423805250036   0.19399834185799544   0.6816135420211479   0.11630289115362488   0.003566006204316518   0.1331358399712277   0.508525772415666   0.5251891559799956   0.7233294585677408   0.828775663514474   0.6559202867000847   0.8619297949407617   0.577525470303529   0.6582184803121754   0.5628943684671404   0.21188388642624228   0.8370945296282681   0.49929189907683397   0.591062212290075   0.8945652708247971   0.4271301147770186   0.9076209208261249   0.80495649751775   0.8208747580387119   0.558487734252015   0.7136225789681294   0.12334295549660218   0.704571866885087   0.5549217280476985   0.5804867389969017   0.6148171830809362   0.17938271090509142   0.8315922694799577   0.7517110754824278   0.9588968963808514   0.3174529159643297   0.25406679917642866   0.09349259517025228   0.39600252791371104   0.10556902953808739
0.4169722695481606   0.5942006960934183   0.804940315623636   0.21100375871329025   0.9898421547711419   0.6865797752672934   0.999983818105886   0.3901290006745783   0.43135442051912687   0.972957196299164   0.8766408626092838   0.6855571337894912   0.8764326924714284   0.39247045730226215   0.26182367952834756   0.5061744228843998   0.0448404229914707   0.6407593818198344   0.30292678314749616   0.1887215069200702   0.790773623815042   0.5472667866495821   0.9069242552337851   0.08315247738198281   0.3738013542668815   0.9530660905561638   0.10198393961014911   0.8721487186686926   0.38395919949573953   0.26648631528887035   0.10200012150426314   0.48201971799411425   0.9526047789766127   0.2935291189897064   0.22535925889497938   0.796462584204623   0.07617208650518427   0.9010586616874443   0.9635355793666318   0.2902881613202231   0.03133166351371356   0.26029927986760987   0.6606087962191356   0.10156665440015294   0.24055803969867154   0.7130324932180278   0.7536845409853505   0.018414177018170125   0.8667566854317901   0.759966402661864   0.6517006013752015   0.14626545834947755   0.48279748593605054   0.49348008737299365   0.5497004798709383   0.6642457403553633   0.5301927069594379   0.19995096838328721   0.3243412209759589   0.8677831561507403   0.4540206204542536   0.29889230669584294   0.36080564160932715   0.5774949948305171
0.42268895694054004   0.038593026828233075   0.7001968453901914   0.47592834043036425   0.18213091724186853   0.3255605336102053   0.9465123044048409   0.4575141634121941   0.31537423181007845   0.5655941309483413   0.2948117030296395   0.31124870506271657   0.832576745874028   0.07211404357534766   0.7451112231587013   0.6470029647073533   0.30238403891459004   0.8721630751920605   0.4207700021827423   0.7792198085566129   0.8483634184603365   0.5732707684962175   0.05996436057341517   0.20172481372609577   0.4256744615197964   0.5346777416679844   0.3597675151832237   0.7257964732957315   0.24354354427792788   0.20911720805777914   0.41325521077838273   0.2682823098835374   0.9281693124678494   0.6435230771094378   0.11844350774874322   0.9570336048208209   0.09559256659382148   0.5714090335340901   0.37333228459004203   0.3100306401134676   0.7932085276792314   0.6992459583420297   0.9525622824072997   0.5308108315568547   0.944845109218895   0.1259751898458122   0.8925979218338845   0.3290860178307589   0.5191706476990986   0.5912974481778278   0.5328304066506608   0.6032895445350274   0.27562710342117075   0.38218024012004864   0.1195751958722781   0.33500723465148996   0.34745779095332135   0.7386571630106108   0.001131688123534872   0.3779736298306691   0.2518652243594999   0.16724812947652065   0.6277994035334928   0.06794298971720152
0.4586566966802684   0.46800217113449094   0.6752371211261932   0.5371321581603469   0.5138115874613735   0.34202698128867876   0.7826391992923086   0.20804614032958793   0.9946409397622747   0.750729533110851   0.2498087926416478   0.6047565957945605   0.719013836341104   0.3685492929908023   0.1302335967693697   0.2697493611430706   0.3715560453877827   0.6298921299801915   0.12910190864583485   0.8917757313124014   0.11969082102828282   0.4626440005036709   0.501302505112342   0.8238327415951999   0.6610341243480145   0.99464182936918   0.8260653839861488   0.28670058343485305   0.147222536886641   0.6526148480805012   0.043426184693840145   0.07865444310526512   0.1525815971243662   0.9018853149696502   0.7936173920521924   0.47389784731070456   0.43356776078326215   0.5333360219788479   0.6633837952828227   0.20414848616763404   0.06201171539547949   0.9034438919986564   0.5342818866369878   0.3123727548552326   0.9423208943671967   0.4407998914949855   0.03297938152464584   0.4885400132600327   0.2812867700191823   0.44615806212580555   0.20691399753849704   0.20183942982517963   0.1340642331325413   0.7935432140453044   0.1634878128446569   0.12318498671991453   0.9814826360081751   0.8916578990756541   0.36987042079246457   0.6492871394092099   0.5479148752249129   0.3583218770968062   0.7064866255096419   0.4451386532415759
0.48590315982943344   0.4548779850981498   0.1722047388726541   0.1327658983863433   0.5435822654622368   0.014078093603164317   0.13922535734800828   0.6442258851263106   0.26229549544305447   0.5679200314773587   0.9323113598095112   0.44238645530113097   0.1282312623105132   0.7743768174320544   0.7688235469648543   0.31920146858121645   0.14674862630233812   0.8827189183564003   0.39895312617238976   0.6699143291720066   0.5988337510774252   0.5243970412595941   0.6924665006627478   0.2247756759304306   0.11293059124799175   0.06951905616144424   0.5202617617900938   0.09200977754408729   0.569348325785755   0.055440962558279926   0.3810364044420855   0.44778389241777666   0.30705283034270053   0.48752093108092115   0.44872504463257423   0.005397437116645731   0.17882156803218732   0.7131441136488668   0.6799014976677199   0.6861959685354293   0.0320729417298492   0.8304251952924665   0.28094837149533014   0.016281639363422796   0.433239190652424   0.3060281540328724   0.5884818708325823   0.7915059634329922   0.32030859940443224   0.23650909787142818   0.06822010904248858   0.6994961858889049   0.7509602736186772   0.18106813531314825   0.6871837046004031   0.2517122934711282   0.44390744327597675   0.693547204232227   0.2384586599678289   0.2463148563544825   0.26508587524378946   0.9804030905833603   0.558557162300109   0.5601188878190532
0.23301293351394023   0.1499778952908938   0.27760879080477885   0.5438372484556304   0.7997737428615163   0.8439497412580214   0.6891269199721965   0.7523312850226382   0.47946514345708396   0.6074406433865932   0.620906810929708   0.052835099133733285   0.7285048698384067   0.42637250807344496   0.9337231063293049   0.8011228056626051   0.2845974265624299   0.7328253038412178   0.695264446361476   0.5548079493081226   0.01951155131864049   0.7524222132578575   0.13670728406136695   0.9946890614890693   0.7864986178047002   0.6024443179669637   0.8590984932565882   0.45085181303343896   0.9867248749431841   0.7584945767089424   0.16997157328439158   0.6985205280108008   0.5072597314861   0.15105393332234915   0.5490647623546836   0.6456854288770675   0.7787548616476934   0.7246814252489042   0.6153416560253788   0.8445626232144624   0.49415743508526344   0.9918561214076864   0.9200772096639028   0.28975467390633985   0.474645883766623   0.23943390814982884   0.7833699256025359   0.2950656124172705   0.6881472659619227   0.636989590182865   0.9242714323459478   0.8442137993838316   0.7014223910187387   0.8784950134739228   0.7542998590615562   0.14569327137303079   0.1941626595326386   0.7274410801515736   0.20523509670687257   0.5000078424959633   0.4154077978849452   0.002759654902669359   0.5898934406814937   0.6554452192815009
0.9212503627996818   0.010903533494982982   0.6698162310175909   0.365690545375161   0.4466044790330588   0.7714696253451542   0.8864463054150551   0.0706249329578905   0.758457213071136   0.13448003516228904   0.9621748730691073   0.22641113357405895   0.057034822052397384   0.2559850216883663   0.20787501400755112   0.0807178622010282   0.8628721625197587   0.5285439415367927   0.0026399173006785553   0.5807100197050649   0.4474643646348136   0.5257842866341234   0.4127464766191848   0.9252648004235641   0.5262140018351319   0.5148807531391404   0.7429302456015938   0.5595742550484031   0.07960952280207308   0.7434111277939862   0.8564839401865387   0.4889493220905125   0.321152309730937   0.6089310926316972   0.8943090671174314   0.26253818851645355   0.26411748767853965   0.35294607094333086   0.6864340531098804   0.18182032631542536   0.40124532515878086   0.8244021294065381   0.6837941358092018   0.6011103066103605   0.9537809605239672   0.2986178427724148   0.271047659190017   0.6758455061867964   0.42756695868883543   0.7837370896332745   0.5281174135884231   0.1162712511383934   0.3479574358867623   0.04032596183928822   0.6716334734018844   0.6273219290478809   0.02680512615582532   0.43139486920759107   0.777324406284453   0.3647837405314273   0.7626876384772857   0.07844879826426016   0.09089035317457267   0.18296341421600196
0.36144231331850485   0.254046668857722   0.4070962173653709   0.5818531076056415   0.4076613527945376   0.9554288260853072   0.1360485581753539   0.9060076014188451   0.9800943941057022   0.17169173645203273   0.6079311445869308   0.7897363502804516   0.6321369582189399   0.1313657746127445   0.9362976711850463   0.1624144212325708   0.6053318320631145   0.6999709054051535   0.15897326490059333   0.7976306807011435   0.8426441935858289   0.6215221071408933   0.06808291172602066   0.6146672664851415   0.48120188026732397   0.3674754382831713   0.6609866943606497   0.03281415887950003   0.0735405274727864   0.41204661219786415   0.5249381361852958   0.12680655746065497   0.09344613336708422   0.2403548757458314   0.9170069915983651   0.3370702071802033   0.4613091751481444   0.1089891011330869   0.9807093204133188   0.1746557859476325   0.8559773430850298   0.40901819572793346   0.8217360555127254   0.377025105246489   0.013333149499201042   0.7874960885870401   0.7536531437867048   0.7623578387613476   0.532131269231877   0.4200206503038688   0.09266644942605506   0.7295436798818474   0.45859074175909065   0.007974038106004696   0.5677283132407592   0.6027371224211925   0.3651446083920064   0.7676191623601732   0.6507213216423942   0.26566691524098923   0.9038354332438621   0.6586300612270863   0.6700120012290753   0.09101112929335671
0.047858090158832155   0.24961186549915296   0.8482759457163499   0.7139860240468677   0.03452494065963111   0.4621157769121128   0.09462280192964503   0.9516281852855202   0.502393671427754   0.042095126608243986   0.0019563525035899637   0.22208450540367272   0.04380292966866341   0.03412108850223929   0.4342280392628307   0.6193473829824803   0.678658321276657   0.266501926142066   0.7835067176204367   0.35368046774149103   0.774822888032795   0.6078718649149796   0.1134947163913613   0.2626693384481343   0.7269647978739628   0.35825999941582665   0.26521877067501143   0.5486833144012666   0.6924398572143317   0.8961442225037138   0.17059596874536642   0.5970551291157464   0.19004618578657764   0.8540490958954698   0.16863961624177645   0.3749706237120737   0.14624325611791422   0.8199280073932306   0.7344115769789457   0.7556232407295934   0.46758493484125724   0.5534260812511645   0.9509048593585091   0.40194277298810244   0.6927620468084623   0.945554216336185   0.8374101429671478   0.13927343453996816   0.9657972489344995   0.5872942169203583   0.5721913722921363   0.5905901201387016   0.27335739172016776   0.6911499944166445   0.4015954035467699   0.9935349910229552   0.08331120593359015   0.8371008985211746   0.2329557873049935   0.6185643673108815   0.9370679498156759   0.01717289112794404   0.4985442103260478   0.862941126581288
0.4694830149744187   0.46374680987677946   0.5476393509675387   0.4609983535931856   0.7767209681659564   0.5181925935405945   0.7102292080003909   0.32172491905321743   0.8109237192314569   0.9308983766202362   0.13803783570825454   0.7311347989145158   0.5375663275112892   0.2397483822035918   0.7364424321614846   0.7375998078915607   0.45425512157769904   0.4026474836824172   0.5034866448564911   0.11903544058067922   0.5171871717620231   0.38547459255447314   0.0049424345304433116   0.2560943139993912   0.04770415678760441   0.9217277826776936   0.4573030835629046   0.7950959604062057   0.270983188621648   0.4035351891370991   0.7470738755625137   0.47337104135298824   0.46005946939019104   0.4726368125168629   0.6090360398542592   0.7422362424384724   0.9224931418789019   0.23288843031327108   0.8725936076927746   0.004636434546911669   0.4682380203012028   0.8302409466308539   0.3691069628362835   0.8856009939662325   0.9510508485391798   0.44476635407638077   0.36416452830584023   0.6295066799668413   0.9033466917515753   0.523038571398687   0.9068614447429356   0.8344107195606356   0.6323635031299273   0.11950338226158795   0.15978756918042186   0.36103967820764743   0.1723040337397363   0.6468665697447251   0.5507515293261627   0.6188034357691751   0.2498108918608344   0.41397813943145395   0.6781579216333881   0.6141670012222634
0.7815728715596316   0.5837371928006001   0.30905095879710454   0.7285660072560309   0.8305220230204519   0.1389708387242193   0.9448864304912643   0.09905932728918966   0.9271753312688765   0.6159322673255322   0.03802498574832872   0.26464860772855403   0.2948118281389492   0.4964288850639443   0.8782374165679069   0.9036089295209067   0.1225077943992129   0.8495623153192192   0.3274858872417442   0.2848054937517316   0.8726969025383785   0.43558417588776527   0.6493279656083562   0.6706384925294683   0.09112403097874691   0.8518469830871652   0.34027700681125167   0.9420724852734373   0.2606020079582951   0.7128761443629459   0.39539057631998736   0.8430131579842477   0.33342667668941856   0.09694387703741364   0.3573655905716586   0.5783645502556936   0.03861484855046936   0.6005149919734694   0.4791281740037518   0.674755620734787   0.9161070541512565   0.7509526766542501   0.15164228676200756   0.38995012698305537   0.043410151612877965   0.31536850076648487   0.5023143211536514   0.7193116344535871   0.9522861206341311   0.46352151767931965   0.1620373143423997   0.7772391491801498   0.691684112675836   0.7506453733163738   0.7666467380224123   0.9342259911959022   0.35825743598641746   0.6537014962789601   0.4092811474507537   0.35586144094020855   0.3196425874359481   0.05318650430549081   0.9301529734470019   0.6811058202054217
0.4035355332846916   0.3022338276512407   0.7785106866849943   0.29115569322236623   0.3601253816718137   0.9868653268847558   0.276196365531343   0.5718440587687791   0.4078392610376826   0.5233438092054362   0.11415905118894332   0.7946049095886293   0.7161551483618466   0.7726984358890624   0.347512313166531   0.8603789183927272   0.35789771237542917   0.11899693961010224   0.9382311657157772   0.5045174774525185   0.038255124939481105   0.06581043530461143   0.008078192268775358   0.823411657247097   0.6347195916547895   0.7635766076533708   0.22956750558378097   0.5322559640247307   0.27459420998297585   0.7767112807686148   0.953371140052438   0.9604119052559515   0.8667549489452933   0.2533674715631787   0.8392120888634946   0.16580699566732227   0.1505998005834466   0.4806690356741163   0.49169977569696366   0.30542807727459514   0.7927020882080175   0.36167209606401407   0.5534686099811864   0.8009105998220766   0.7544469632685363   0.2958616607594026   0.545390417712411   0.9774989425749797   0.11972737161374684   0.5322850531060319   0.31582291212863006   0.44524297855024897   0.845133161630771   0.7555737723374171   0.36245177207619206   0.4848310732942974   0.9783782126854778   0.5022063007742383   0.5232396832126974   0.31902407762697516   0.8277784121020312   0.021537265100122015   0.031539907515733774   0.01359600035237998
0.03507632389401375   0.6598651690361079   0.4780712975345474   0.21268540053030338   0.28062936062547744   0.3640035082767053   0.9326808798221363   0.23518645795532372   0.16090198901173058   0.8317184551706734   0.6168579676935063   0.7899434794050747   0.31576882738095957   0.0761446828332564   0.25440619561731426   0.30511240611077733   0.33739061469548176   0.573938382059018   0.7311665124046168   0.9860883284838022   0.5096122025934506   0.552401116958896   0.6996266048888831   0.9724923281314223   0.47453587869943686   0.8925359479227881   0.22155530735433565   0.7598069276011189   0.19390651807395942   0.5285324396460828   0.2888744275321993   0.5246204696457951   0.03300452906222885   0.6968139844754094   0.672016459838693   0.7346769902407204   0.7172357016812693   0.620669301642153   0.4176102642213787   0.42956458412994303   0.3798450869857875   0.04673091958313491   0.6864437518167619   0.44347625564614085   0.8702328843923369   0.49432980262423887   0.9868171469278788   0.4709839275147186   0.3956970056929   0.6017938547014507   0.7652618395735432   0.7111769999135997   0.20179048761894058   0.07326141505536794   0.4763874120413439   0.18655653026780464   0.16878595855671175   0.37644743057995855   0.804370952202651   0.45187954002708425   0.4515502568754425   0.7557781289378056   0.3867606879812723   0.02231495589714119
0.07170516988965497   0.7090472093546707   0.7003169361645104   0.5788387002510004   0.20147228549731808   0.21471740673043183   0.7134997892366316   0.10785477273628172   0.8057752798044181   0.6129235520289811   0.9482379496630884   0.39667777282268196   0.6039847921854775   0.5396621369736131   0.4718505376217445   0.21012124255487732   0.4351988336287657   0.1632147063936546   0.6674795854190936   0.7582417025277931   0.9836485767533233   0.407436577455849   0.2807188974378213   0.7359267466306518   0.9119434068636683   0.6983893681011784   0.5804019612733109   0.15708804637965154   0.7104711213663502   0.48367196137074653   0.8669021720366794   0.049233273643369824   0.9046958415619322   0.8707484093417655   0.9186642223735909   0.6525555008206879   0.30071104937645465   0.3310862723681523   0.4468136847518464   0.44243425826581056   0.865512215747689   0.1678715659744977   0.7793340993327529   0.6841925557380175   0.8818636389943657   0.7604349885186487   0.4986152018949315   0.9482658091073656   0.9699202321306974   0.06204562041747035   0.9182132406216206   0.7911777627277141   0.25944911076434723   0.5783736590467238   0.05131106858494123   0.7419444890843443   0.3547532692024151   0.7076252497049583   0.13264684621135028   0.08938898826365638   0.054042219825960455   0.3765389773368061   0.6858331614595039   0.6469547299978459
0.1885300040782715   0.20866741136230837   0.906499062126751   0.9627621742598284   0.3066663650839058   0.44823242284365966   0.4078838602318195   0.014496365152462711   0.3367461329532084   0.3861868024261893   0.4896706196101989   0.22331860242474863   0.07729702218886111   0.8078131433794655   0.4383595510252577   0.48137411334040436   0.722543752986446   0.10018789367450712   0.3057127048139074   0.391985125076748   0.6685015331604856   0.723648916337701   0.6198795433544035   0.7450303950789022   0.479971529082214   0.5149815049753926   0.7133804812276525   0.7822682208190739   0.17330516399830825   0.06674908213173301   0.305496620995833   0.7677718556666112   0.8365590310450999   0.6805622797055437   0.8158260013856341   0.5444532532418626   0.7592620088562387   0.8727491363260782   0.3774664503603764   0.06307913990145814   0.03671825586979277   0.7725612426515711   0.07175374554646902   0.6710940148247101   0.3682167227093072   0.04891232631387004   0.4518742021920655   0.926063619745808   0.8882451936270932   0.5339308213384774   0.7384937209644129   0.14379539892673407   0.714940029628785   0.46718173920674433   0.43299709996857993   0.3760235432601229   0.8783809985836851   0.7866194595012007   0.6171710985829458   0.8315702900182603   0.11911898972744632   0.9138703231751225   0.23970464822256937   0.7684911501168022
0.08240073385765355   0.14130908052355137   0.16795090267610038   0.09739713529209212   0.7141840111483463   0.09239675420968134   0.7160767004840349   0.1713335155462842   0.8259388175212531   0.5584659328712039   0.9775829795196219   0.02753811661955014   0.11099878789246816   0.09128419366445961   0.5445858795510421   0.6515145733594272   0.23261778930878307   0.30466473416325895   0.9274147809680963   0.8199442833411669   0.11349879958133677   0.3907944109881365   0.6877101327455268   0.051453133224364615   0.031098065723683222   0.24948533046458513   0.5197592300694265   0.9540559979322725   0.3169140545753369   0.15708857625490377   0.8036825295853915   0.7827224823859883   0.4909752370540838   0.5986226433836999   0.8260995500657696   0.7551843657664381   0.37997644916161566   0.5073384497192402   0.28151367051472753   0.1036697924070109   0.14735865985283256   0.20267371555598127   0.35409888954663127   0.28372550906584404   0.0338598602714958   0.8118793045678447   0.6663887568011044   0.23227237584147942   0.002761794547812572   0.5623939741032596   0.1466295267316779   0.27821637790920695   0.6858477399724756   0.40530539784835584   0.3429469971462863   0.49549389552321865   0.19487250291839187   0.8066827544646561   0.5168474470805167   0.7403095297567805   0.8148960537567762   0.29934430474541585   0.23533377656578913   0.6366397373497696
0.6675373939039436   0.0966705891894346   0.8812348870191579   0.35291422828392555   0.6336775336324478   0.2847912846215898   0.21484613021805343   0.12064185244244614   0.6309157390846353   0.7223973105183302   0.06821660348637551   0.8424254745332392   0.9450679991121597   0.31709191266997433   0.7252696063400892   0.3469315790100206   0.7501954961937678   0.5104091582053183   0.20842215925957253   0.60662204925324   0.9352994424369916   0.21106485345990242   0.9730883826937834   0.9699823119034705   0.26776204853304786   0.11439426427046782   0.09185349567462556   0.6170680836195449   0.6340845149006   0.829602979648878   0.8770073654565721   0.4964262311770988   0.0031687758159646973   0.10720566913054783   0.8087907619701966   0.6540007566438596   0.058100776703805056   0.7901137564605735   0.08352115563010742   0.307069177633839   0.3079052805100373   0.27970459825525523   0.8750989963705349   0.7004471283805989   0.3726058380730457   0.06863974479535283   0.9020106136767515   0.7304648164771285   0.10484378953999784   0.954245480524885   0.810157118002126   0.11339673285758355   0.4707592746393979   0.12464250087600699   0.9331497525455538   0.6169705016804848   0.4675904988234332   0.017436831745459166   0.12435899057535718   0.9629697450366252   0.4094897221196281   0.22732307528488566   0.040837834945249764   0.6559005674027862
0.10158444160959082   0.9476184770296304   0.16573883857471486   0.9554534390221874   0.7289786035365451   0.8789787322342776   0.2637282248979634   0.2249886225450589   0.6241348139965472   0.9247332517093926   0.4535711068958374   0.11159188968747534   0.1533755393571494   0.8000907508333857   0.5204213543502836   0.49462138800699057   0.6857850405337163   0.7826539190879265   0.39606236377492643   0.5316516429703653   0.27629531841408816   0.5553308438030408   0.35522452882967664   0.875751075567579   0.17471087680449732   0.6077123667734103   0.18948569025496179   0.9202976365453918   0.44573227326795223   0.7287336345391328   0.9257574653569984   0.6953090140003328   0.821597459271405   0.8040003828297402   0.472186358461161   0.5837171243128575   0.6682219199142556   0.003909631996354563   0.9517650041108774   0.08909573630586694   0.9824368793805394   0.2212557129084281   0.555702640335951   0.5574440933355016   0.7061415609664512   0.6659248691053873   0.20047811150627434   0.6816930177679226   0.5314306841619539   0.058212502331976945   0.010992421251312565   0.7613953812225308   0.08569841089400168   0.3294788677928442   0.08523495589431414   0.06608636722219799   0.26410095162259667   0.525478484963104   0.6130485974331531   0.4823692429093405   0.5958790317083411   0.5215688529667494   0.6612835933222757   0.39327350660347354
0.6134421523278017   0.3003131400583213   0.10558095298632472   0.835829413267972   0.9073005913613504   0.6343882709529339   0.9051028414800504   0.1541363955000494   0.37586990719939656   0.576175768620957   0.8941104202287378   0.39274101427751856   0.2901714963053949   0.24669690082811288   0.8088754643344237   0.3266546470553206   0.026070544682798204   0.7212184158650089   0.19582686690127055   0.8442854041459801   0.4301915129744571   0.19964956289825947   0.5345432735789948   0.45101189754250653   0.8167493606466554   0.8993364228399382   0.4289623205926701   0.6151824842745346   0.9094487692853049   0.26494815188700416   0.5238594791126198   0.46104608877448516   0.5335788620859084   0.6887723832660472   0.6297490588838819   0.0683050744969666   0.2434073657805135   0.44207548243793426   0.8208735945494582   0.741650427441646   0.2173368210977153   0.7208570665729254   0.6250467276481877   0.8973650232956659   0.7871453081232581   0.521207503674666   0.09050345406919286   0.4463531257531594   0.9703959474766027   0.6218710808347278   0.6615411334765228   0.8311706414786247   0.06094717819129779   0.3569229289477236   0.13768165436390306   0.37012455270413963   0.5273683161053894   0.6681505456816764   0.5079325954800211   0.30181947820717303   0.2839609503248759   0.22607506324374219   0.6870590009305629   0.560169050765527
0.0666241292271606   0.5052179966708168   0.062012273282375276   0.6628040274698611   0.27947882110390243   0.984010492996151   0.9715088192131824   0.21645090171670173   0.3090828736272997   0.36213941216142315   0.30996768573665967   0.38528026023807693   0.2481356954360019   0.005216483213699588   0.1722860313727566   0.015155707533937322   0.7207673793306125   0.33706593753202313   0.6643534358927354   0.7133362293267643   0.43680642900573663   0.11099087428828097   0.9772944349621725   0.1531671785612373   0.37018229977857603   0.6057728776174641   0.9152821616797973   0.4903631510913762   0.0907034786746736   0.6217623846213133   0.9437733424666148   0.27391224937467445   0.7816206050473739   0.2596229724598901   0.6338056567299551   0.8886319891365976   0.533484909611372   0.2544064892461905   0.46151962535719854   0.8734762816026602   0.8127175302807595   0.9173405517141674   0.797166189464463   0.16014005227589592   0.37591110127502286   0.8063496774258864   0.8198717545022907   0.006972873714658609   0.0057288014964468545   0.20057679980842222   0.9045895928224934   0.5166097226232824   0.9150253228217733   0.578814415187109   0.9608162503558786   0.24269747324860794   0.13340471777439936   0.3191914427272189   0.3270105936259235   0.3540654841120104   0.5999198081630274   0.06478495348102839   0.865490968268725   0.48058920250935017
0.7872022778822678   0.14744440176686105   0.06832477880426184   0.32044915023345427   0.41129117660724496   0.34109472434097465   0.24845302430197122   0.31347627651879567   0.4055623751107981   0.1405179245325524   0.34386343147947784   0.7968665538955132   0.4905370522890249   0.5617035093454434   0.38304718112359926   0.5541690806469053   0.3571323345146255   0.24251206661822455   0.05603658749767576   0.20010359653489493   0.7572125263515982   0.17772711313719616   0.19054561922895083   0.7195143940255447   0.9700102484693303   0.03028271137033512   0.12222084042468898   0.39906524379209046   0.5587190718620854   0.6891879870293605   0.8737678161227177   0.08558896727329483   0.1531566967512872   0.548670062496808   0.52990438464324   0.2887224133777816   0.6626196444622623   0.9869665531513646   0.14685720351964068   0.7345533327308763   0.30548730994763684   0.7444544865331401   0.09082061602196492   0.5344497361959814   0.5482747835960387   0.5667273733959439   0.9002749967930141   0.8149353421704366   0.5782645351267084   0.5364446620256088   0.7780541563683251   0.41587009837834615   0.019545463264623027   0.8472566749962483   0.9042863402456074   0.3302811311050513   0.8663887665133359   0.29858661249944024   0.3743819556023675   0.04155871772726972   0.2037691220510735   0.31162005934807563   0.22752475208272677   0.30700538499639346
0.8982818121034367   0.5671655728149356   0.13670413606076184   0.772555648800412   0.350007028507398   0.00043819941899169703   0.23642913926774775   0.9576203066299754   0.7717424933806897   0.4639935373933829   0.45837498289942263   0.5417502082516293   0.7521970301160666   0.6167368623971347   0.5540886426538153   0.21146907714657803   0.8858082636027308   0.31815024989769436   0.1797066870514478   0.16991035941930832   0.6820391415516573   0.00653019054961869   0.952181934968721   0.8629049744229149   0.7837573294482206   0.4393646177346831   0.8154777989079591   0.09034932562250278   0.4337503009408226   0.4389264183156914   0.5790486596402115   0.13272901899252731   0.6620078075601329   0.9749328809223085   0.12067367674078881   0.590978810740898   0.9098107774440662   0.35819601852517385   0.5665850340869736   0.37950973359431994   0.02400251384133543   0.04004576862747952   0.38687834703552576   0.20959937417501162   0.3419633722896781   0.03351557807786083   0.4346964120668047   0.34669439975209676   0.5582060428414575   0.5941509603431777   0.6192186131588455   0.25634507412959395   0.12445574190063487   0.15522454202748634   0.040169953518634116   0.12361605513706667   0.46244793434050196   0.18029166110517786   0.9194962767778453   0.5326372443961687   0.5526371568964357   0.822095642580004   0.35291124269087176   0.15312751080184875
0.5286346430551002   0.7820498739525245   0.966032895655346   0.9435281366268371   0.18667127076542217   0.7485342958746637   0.5313364835885412   0.5968337368747404   0.6284652279239646   0.1543833355314859   0.9121178704296957   0.3404886627451464   0.5040094860233298   0.9991587935039995   0.8719479169110617   0.21687260760807972   0.041561551682827866   0.8188671323988217   0.9524516401332163   0.684235363211911   0.48892439478639216   0.9967714898188177   0.5995403974423446   0.5311078524100623   0.9602897517312919   0.2147216158662932   0.6335075017869986   0.5875797157832252   0.7736184809658697   0.4661873199916296   0.10217101819845725   0.9907459789084848   0.14515325304190507   0.3118039844601437   0.19005314776876153   0.6502573161633385   0.6411437670185752   0.3126451909561441   0.3181052308576999   0.43338470855525874   0.5995822153357474   0.49377805855732243   0.3656535907244836   0.7491493453433478   0.1106578205493552   0.4970065687385048   0.7661131932821391   0.21804149293328542   0.1503680688180633   0.28228495287221156   0.13260569149514057   0.6304617771500602   0.37674958785219353   0.816097632880582   0.030434673296683312   0.6397157982415754   0.23159633481028846   0.5042936484204383   0.8403815255279218   0.989458482078237   0.5904525677917132   0.19164845746429418   0.5222762946702219   0.5560737735229782
0.9908703524559659   0.6978703989069718   0.15662270394573824   0.8069244281796305   0.8802125319066106   0.20086383016846696   0.3905095106635992   0.588882935246345   0.7298444630885473   0.9185788772962554   0.2579038191684586   0.9584211580962848   0.3530948752363538   0.10248124441567341   0.2274691458717753   0.31870535985470944   0.12149854042606534   0.5981875959952351   0.3870876203438535   0.3292468777764725   0.5310459726343522   0.4065391385309409   0.8648113256736316   0.7731731042534943   0.5401756201783863   0.7086687396239693   0.7081886217278934   0.9662486760738638   0.6599630882717756   0.5078049094555023   0.3176791110642942   0.3773657408275188   0.9301186251832283   0.5892260321592468   0.05977529189583561   0.4189445827312339   0.5770237499468744   0.48674478774357344   0.8323061460240603   0.10023922287652451   0.45552520952080916   0.8885571917483384   0.4452185256802068   0.770992345100052   0.9244792368864571   0.4820180532173974   0.5804072000065752   0.9978192408465577   0.3843036167080708   0.7733493135934282   0.8722185782786818   0.03157056477269393   0.7243405284362952   0.26554440413792596   0.5545394672143876   0.6542048239451752   0.7942219032530669   0.6763183719786791   0.494764175318552   0.23526024121394123   0.21719815330619233   0.18957358423510565   0.6624580292944917   0.13502101833741673
0.7616729437853832   0.3010163924867673   0.21723950361428485   0.3640286732373647   0.8371937068989261   0.8189983392693699   0.6368323036077097   0.36620943239080694   0.4528900901908554   0.04564902567594172   0.7646137253290278   0.334638867618113   0.7285495617545603   0.7801046215380157   0.21007425811464028   0.6804340436729378   0.9343276585014935   0.10378624955933669   0.7153100827960883   0.4451738024589966   0.7171295051953012   0.9142126653242311   0.05285205350159662   0.31015278412157987   0.955456561409918   0.6131962728374637   0.8356125498873118   0.9461241108842152   0.11826285451099178   0.7941979335680938   0.19878024627960209   0.5799146784934083   0.6653727643201364   0.748548907892152   0.43416652095057423   0.24527581087529524   0.936823202565576   0.9684442863541363   0.22409226283593395   0.5648417672023573   0.0024955440640826248   0.8646580367947996   0.5087821800398457   0.11966796474336078   0.2853660388687815   0.9504453714705686   0.45593012653824905   0.8095151806217808   0.32990947745886356   0.33724909863310487   0.6203175766509372   0.8633910697375657   0.2116466229478718   0.543051165065011   0.4215373303713352   0.28347639124415747   0.5462738586277354   0.794502257172859   0.9873708094207609   0.03820058036886221   0.6094506560621593   0.8260579708187228   0.763278546584827   0.4733588131665048
0.6069551119980767   0.9613999340239231   0.2544963665449813   0.353690848423144   0.3215890731292952   0.010954562553354573   0.7985662400067323   0.5441756678013632   0.9916795956704316   0.6737054639202497   0.178248663355795   0.6807845980637974   0.7800329727225599   0.1306542988552386   0.7567113329844598   0.39730820681964   0.23375911409482442   0.3361520416823796   0.7693405235636989   0.3591076264507778   0.6243084580326651   0.5100940708636569   0.006061976978871923   0.885748813284273   0.01735334603458839   0.5486941368397337   0.7515656104338906   0.532057964861129   0.6957642729052932   0.5377395742863791   0.9529993704271583   0.9878822970597658   0.7040846772348616   0.8640341103661294   0.7747507070713633   0.30709769899596834   0.9240517045123017   0.7333798115108908   0.018039374086903447   0.9097894921763283   0.6902925904174773   0.3972277698285112   0.24869885052320453   0.5506818657255506   0.06598413238481217   0.8871336989648544   0.2426368735443326   0.6649330524412775   0.048630786350223776   0.33843956212512066   0.491071263110442   0.1328750875801486   0.3528665134449306   0.8006999878387415   0.5380718926832837   0.1449927905203828   0.648781836210069   0.9366658774726121   0.7633211856119204   0.8378950915244144   0.7247301316977673   0.2032860659617213   0.7452818115250169   0.9281055993480861
0.034437541280290085   0.8060582961332101   0.49658296100181243   0.3774237336225356   0.9684534088954779   0.9189245971683557   0.2539460874574798   0.712490681181258   0.9198226225452542   0.580485035043235   0.7628748243470378   0.5796155936011095   0.5669561091003236   0.7797850472044935   0.2248029316637541   0.43462280308072665   0.9181742728902546   0.8431191697318814   0.4614817460518337   0.5967277115563122   0.19344414119248715   0.6398331037701601   0.7161999345268167   0.6686221122082261   0.15900659991219707   0.83377480763695   0.2196169735250043   0.2911983785856905   0.19055319101671916   0.9148502104685943   0.9656708860675245   0.5787076974044324   0.27073056847146504   0.3343651754253592   0.20279606172048673   0.9990921038033229   0.7037744593711415   0.5545801282208657   0.9779931300567326   0.5644693007225963   0.7856001864808869   0.7114609584889843   0.5165113840048989   0.9677415891662842   0.5921560452883998   0.07162785471882421   0.8003114494780822   0.2991194769580581   0.43314944537620276   0.2378530470818742   0.5806944759530779   0.007921098372367628   0.2425962543594836   0.32300283661327994   0.6150235898855534   0.4292134009679352   0.9718656858880186   0.9886376611879207   0.4122275281650667   0.4301212971646123   0.2680912265168771   0.43405753296705507   0.43423439810833403   0.865651996442016
0.48249104003599014   0.7225965744780708   0.9177230141034352   0.8979104072757318   0.8903349947475904   0.6509687197592465   0.1174115646253529   0.5987909303176737   0.45718554937138756   0.4131156726773723   0.536717088672275   0.5908698319453061   0.21458929501190396   0.09011283606409237   0.9216934987867216   0.16165643097737087   0.24272360912388538   0.10147517487617162   0.5094659706216549   0.7315351338127586   0.9746323826070082   0.6674176419091166   0.07523157251332085   0.8658831373707426   0.4921413425710181   0.9448210674310458   0.15750855840988573   0.9679727300950108   0.6018063478234278   0.29385234767179924   0.04009699378453284   0.36918179977733717   0.1446207984520402   0.8807366749944269   0.5033799051122578   0.778311967832031   0.9300315034401363   0.7906238389303345   0.5816864063255363   0.6166555368546602   0.6873078943162508   0.6891486640541629   0.07222043570388134   0.8851204030419016   0.7126755117092426   0.021731022145046328   0.9969888631905605   0.019237265671158934   0.22053416913822446   0.07690995471400054   0.8394803047806747   0.05126453557614807   0.6187278213147966   0.7830576070422013   0.7993833109961419   0.682082735798811   0.47410702286275647   0.9023209320477744   0.2960034058838841   0.9037707679667798   0.5440755194226202   0.1116970931174399   0.7143169995583478   0.2871152311121196
0.8567676251063694   0.422548429063277   0.6420965638544665   0.401994828070218   0.14409211339712677   0.4008174069182307   0.645107700663906   0.3827575623990591   0.9235579442589023   0.3239074522042302   0.8056273958832313   0.33149302682291104   0.3048301229441056   0.5408498451620288   0.006244084887089343   0.6494102910241001   0.8307231000813492   0.6385289131142544   0.7102406790032053   0.7456395230573203   0.2866475806587289   0.5268318199968145   0.9959236794448575   0.45852429194520067   0.4298799555523596   0.1042833909335375   0.353827115590391   0.05652946387498263   0.28578784215523284   0.7034659840153068   0.708719414926485   0.6737719014759236   0.36222989789633053   0.3795585318110767   0.9030920190432538   0.3422788746530125   0.05739977495222493   0.8387086866490479   0.8968479341561644   0.6928685836289123   0.22667667487087578   0.2001797735347934   0.18660725515295915   0.9472290605715921   0.9400290942121469   0.6733479535379789   0.19068357570810165   0.48870476862639145   0.5101491386597873   0.5690645626044414   0.8368564601177106   0.4321753047514088   0.22436129650455444   0.8655985785891346   0.12813704519122565   0.7584034032754853   0.862131398608224   0.4860400467780579   0.22504502614797187   0.41612452862247273   0.804731623655999   0.64733136012901   0.32819709199180747   0.7232559449935604
0.5780549487851232   0.44715158659421667   0.14158983683884832   0.7760268844219683   0.6380258545729763   0.7738036330562378   0.9509062611307466   0.28732211579557687   0.12787671591318908   0.2047390704517964   0.114049801013036   0.855146811044168   0.9035154194086347   0.3391404918626618   0.9859127558218104   0.0967434077686828   0.041384020800410704   0.8531004450846039   0.7608677296738384   0.68061887914621   0.23665239714441172   0.20576908495559382   0.432670637682031   0.9573629341526496   0.6585974483592885   0.7586174983613772   0.2910808008431827   0.18133604973068135   0.020571593786312167   0.9848138653051393   0.34017453971243605   0.8940139339351045   0.8926948778731231   0.7800747948533429   0.22612473869940006   0.03886712289093644   0.9891794584644885   0.4409343029906811   0.24021198287758969   0.9421237151222537   0.9477954376640778   0.5878338579060771   0.47934425320375124   0.2615048359760436   0.711143040519666   0.38206477295048336   0.0466736155217202   0.30414190182339396   0.05254559216037754   0.6234472745891062   0.7555928146785374   0.1228058520927126   0.03197399837406538   0.638633409283967   0.41541827496610145   0.2287919181576081   0.1392791205009423   0.858558614430624   0.1892935362667014   0.18992479526667166   0.1500996620364538   0.41762431143994294   0.9490815533891117   0.247801080144418
0.20230422437237602   0.8297904535338658   0.4697373001853605   0.9862962441683744   0.49116118385270996   0.4477256805833824   0.42306368466364025   0.6821543423449804   0.43861559169233244   0.8242784059942762   0.6674708699851027   0.5593484902522678   0.40664159331826705   0.18564499671030926   0.2520525950190013   0.3305565720946598   0.2673624728173248   0.32708638227968523   0.06275905875229991   0.14063177682798808   0.11726281078087097   0.9094620708397423   0.1136775053631882   0.8928306966835701   0.9149585864084949   0.0796716173058765   0.6439402051778277   0.9065344525151957   0.42379740255578496   0.6319459367224941   0.22087652051418746   0.22438011017021522   0.9851818108634525   0.8076675307282178   0.5534056505290846   0.6650316199179473   0.5785402175451855   0.6220225340179086   0.30135305551008335   0.33447504782328763   0.3111777447278607   0.2949361517382234   0.23859399675778345   0.19384327099529955   0.19391493394698972   0.3854740808984811   0.12491649139459524   0.30101257431172945   0.2789563475384948   0.3058024635926046   0.4809762862167675   0.3944781217965338   0.8551589449827098   0.6738565268701106   0.2600997657025801   0.17009801162631857   0.8699771341192573   0.8661889961418926   0.7066941151734953   0.5050663917083712   0.29143691657407184   0.24416646212398402   0.40534105966341205   0.17059134388508357
0.9802591718462111   0.9492303103857607   0.16674706290562857   0.976748072889784   0.7863442378992215   0.5637562294872795   0.04183057151103334   0.6757354985780546   0.5073878903607266   0.2579537658946749   0.5608542852942658   0.2812573767815208   0.6522289453780168   0.5840972390245643   0.30075451959168575   0.1111593651552022   0.7822518112587595   0.7179082428826717   0.5940604044181904   0.606092973446831   0.4908148946846877   0.47374178075868767   0.18871934475477833   0.4355016295617474   0.5105557228384765   0.5245114703729271   0.021972281849149757   0.4587535566719634   0.7242114849392551   0.9607552408856476   0.9801417103381164   0.7830180580939088   0.21682359457852846   0.7028014749909727   0.4192874250438506   0.501760681312388   0.5645946492005116   0.11870423596640828   0.11853290545216484   0.3906013161571858   0.7823428379417521   0.40079599308373653   0.5244725010339745   0.7845083427103549   0.2915279432570644   0.9270542123250489   0.33575315627919616   0.34900671314860743   0.7809722204185878   0.4025427419521218   0.3137808744300464   0.890253156476644   0.05676073547933273   0.44178750106647424   0.33363916409192995   0.10723509838273527   0.8399371409008043   0.7389860260755016   0.9143517390480794   0.6054744170703472   0.2753424917002927   0.6202817901090933   0.7958188335959145   0.21487310091316142
0.4929996537585406   0.21948579702535675   0.27134633256194   0.4303647582028066   0.20147171050147622   0.2924315847003079   0.9355931762827439   0.08135804505419918   0.4204994900828884   0.8898888427481861   0.6218123018526975   0.19110488857755512   0.36373875460355565   0.44810134168171184   0.28817313776076753   0.08386979019481984   0.5238016137027514   0.7091153156062102   0.37382139871268816   0.4783953731244726   0.24845912200245868   0.08883352549711691   0.5780025651167736   0.26352227221131114   0.7554594682439181   0.8693477284717601   0.3066562325548336   0.8331575140085046   0.5539877577424419   0.5769161437714523   0.3710630562720897   0.7517994689543054   0.13348826765955352   0.6870273010232661   0.7492507544193922   0.5606945803767502   0.7697495130559979   0.2389259593415543   0.4610776166586247   0.4768247901819304   0.24594789935324654   0.529810643735344   0.0872562179459365   0.9984294170574578   0.9974887773507879   0.44097711823822716   0.5092536528291629   0.7349071448461467   0.24202930910686973   0.5716293897664669   0.20259742027432928   0.9017496308376421   0.6880415513644279   0.9947132459950148   0.8315343640022396   0.14995016188333674   0.5545532837048743   0.3076859449717486   0.0822836095828474   0.5892555815065864   0.7848037706488764   0.0687599856301943   0.6212059929242227   0.11243079132465601
0.53885587129563   0.5389493418948502   0.5339497749782862   0.11400137426719816   0.5413670939448421   0.0979722236566231   0.02469612214912334   0.3790942294210515   0.2993377848379723   0.5263428338901561   0.8220987018747941   0.47734459858340933   0.6112962334735444   0.5316295878951414   0.9905643378725545   0.3273944367000726   0.056742949768670135   0.22394364292339278   0.9082807282897071   0.7381388551934862   0.2719391791197937   0.1551836572931985   0.28707473536548433   0.6257080638688302   0.7330833078241638   0.6162343153983483   0.7531249603871981   0.511706689601632   0.19171621387932172   0.5182620917417251   0.7284288382380748   0.13261246018058054   0.8923784290413495   0.9919192578515691   0.9063301363632807   0.6552678615971712   0.28108219556780495   0.46028966995642767   0.9157657984907263   0.3278734248970986   0.2243392457991348   0.2363460270330349   0.0074850702010191995   0.5897345697036124   0.9524000666793411   0.0811623697398364   0.7204103348355348   0.9640265058347822   0.21931675885517732   0.46492805434148815   0.9672853744483367   0.45231981623315026   0.027600544975855606   0.946665962599763   0.23885653621026198   0.3197073560525697   0.1352221159345062   0.9547467047481939   0.3325263998469813   0.6644394944553985   0.8541399203667013   0.4944570347917663   0.41676060135625503   0.3365660695583
0.6298006745675665   0.25811100775873136   0.4092755311552358   0.7468314998546876   0.6774006078882254   0.17694863801889496   0.6888651963197009   0.7828049940199053   0.45808384903304805   0.7120205836774068   0.7215798218713642   0.330485177786755   0.43048330405719243   0.7653546210776438   0.4827232856611022   0.010777821734185301   0.29526118812268626   0.8106079163294498   0.1501968858141209   0.3463383272787868   0.441121267755985   0.3161508815376836   0.7334362844578659   0.009772257720486767   0.8113205931884184   0.05803987377895225   0.3241607533026301   0.2629407578657992   0.1339199853001931   0.8810912357600573   0.6352955569829292   0.4801357638458939   0.675836136267145   0.16907065208265046   0.913715735111565   0.14965058605913886   0.2453528322099526   0.40371603100500664   0.4309924494504628   0.13887276432495355   0.9500916440872664   0.5931081146755567   0.28079556363634184   0.7925344370461668   0.5089703763312814   0.2769572331378731   0.5473592791784759   0.78276217932568   0.697649783142863   0.21891735935892087   0.22319852587584585   0.5198214214598809   0.5637297978426699   0.3378261235988636   0.5879029688929167   0.039685657613986944   0.8878936615755247   0.16875547151621315   0.6741872337813517   0.8900350715548481   0.6425408293655722   0.7650394405112065   0.24319478433088892   0.7511623072298945
0.6924491852783058   0.17193132583564977   0.9623992206945471   0.9586278701837277   0.1834788089470244   0.8949740926977766   0.4150399415160711   0.1758656908580477   0.48582902580416143   0.6760567333388557   0.19184141564022528   0.6560442693981668   0.9220992279614916   0.3382306097399922   0.6039384467473086   0.6163586117841799   0.03420556638596683   0.16947513822377905   0.9297512129659569   0.7263235402293319   0.39166473702039467   0.40443569771257254   0.6865564286350679   0.9751612329994372   0.6992155517420888   0.23250437187692274   0.724157207940521   0.01653336281570955   0.5157367427950644   0.3375302791791461   0.3091172664244498   0.8406676719576619   0.02990771699090302   0.6614735458402903   0.11727585078422456   0.184623402559495   0.10780848902941141   0.32324293610029814   0.513337404036916   0.5682647907753151   0.07360292264344459   0.15376779787651912   0.5835861910709591   0.8419412505459832   0.68193818562305   0.7493321001639466   0.897029762435891   0.866780017546546   0.982722633880961   0.5168277282870238   0.17287255449537017   0.8502466547308364   0.4669858910858966   0.17929744910787773   0.8637552880709204   0.009578982773174562   0.4370781740949936   0.5178239032675874   0.7464794372866957   0.8249555802136795   0.3292696850655822   0.19458096716728926   0.23314203324977983   0.2566907894383645
0.2556667624221376   0.04081316929077016   0.6495558421788208   0.41474953889238125   0.5737285767990876   0.2914810691268236   0.7525260797429296   0.5479695213458353   0.5910059429181266   0.7746533408397998   0.5796535252475594   0.6977228666149988   0.12402005183222997   0.595355891731922   0.7158982371766391   0.6881438838418243   0.6869418777372364   0.0775319884643346   0.9694187998899433   0.8631883036281447   0.3576721926716542   0.8829510212970453   0.7362767666401635   0.6064975141897803   0.10200543024951658   0.8421378520062751   0.08672092446134275   0.19174797529739898   0.528276853450429   0.5506567828794516   0.3341948447184131   0.6437784539515637   0.9372709105323024   0.7760034420396519   0.7545413194708537   0.9460555873365648   0.8132508587000724   0.18064755030772983   0.03864308229421452   0.2579117034947406   0.126308980962836   0.10311556184339525   0.06922428240427121   0.3947233998665958   0.7686367882911819   0.22016454054634993   0.3329475157641077   0.7882258856768156   0.6666313580416652   0.37802668854007476   0.24622659130276497   0.5964779103794167   0.1383545045912363   0.8273699056606232   0.9120317465843518   0.9526994564278529   0.20108359405893397   0.05136646362097132   0.15749042711349823   0.006643869091288029   0.3878327353588616   0.8707189133132415   0.11884734481928372   0.7487321655965474
0.2615237543960256   0.7676033514698463   0.049623062415012506   0.3540087657299516   0.4928869661048438   0.5474388109234963   0.7166755466509048   0.565782880053136   0.8262556080631785   0.16941212238342154   0.4704489553481398   0.9693049696737194   0.6879011034719422   0.3420422167227984   0.558417208763788   0.016605513245866517   0.4868175094130083   0.2906757531018271   0.4009267816502897   0.009961644154578488   0.09898477405414666   0.4199568397885856   0.282079436831006   0.261229478558031   0.837461019658121   0.6523534883187394   0.23245637441599348   0.9072207128280794   0.3445740535532773   0.10491467739524306   0.5157808277650887   0.3414378327749434   0.5183184454900988   0.9355025550118216   0.045331872416948894   0.37213286310122395   0.8304173420181565   0.5934603382890231   0.48691466365316094   0.35552734985535744   0.3435998326051482   0.30278458518719603   0.08598788200287125   0.345565705700779   0.24461505855100157   0.8828277453986104   0.8039084451718652   0.08433622714274794   0.4071540388928805   0.23047425707987107   0.5714520707558718   0.17711551431466854   0.06257998533960324   0.125559579684628   0.055671242990783056   0.8356776815397252   0.5442615398495045   0.1900570246728065   0.010339370573834165   0.4635448184385012   0.713844197831348   0.5965966863837834   0.5234247069206732   0.10801746858314375
0.3702443652261998   0.29381210119658735   0.43743682491780195   0.7624517628823648   0.12562930667519823   0.41098435579797693   0.6335283797459367   0.6781155357396168   0.7184752677823177   0.18051009871810583   0.06207630899006495   0.5010000214249483   0.6558952824427144   0.054950519033477835   0.0064050659992818905   0.6653223398852232   0.11163374259320996   0.8648934943606713   0.9960656954254478   0.20177752144672192   0.39778954476186196   0.26829680797688793   0.4726409885047745   0.09376005286357818   0.02754517953566215   0.9744847067803006   0.035204163586972544   0.3313082899812134   0.9019158728604639   0.5635003509823237   0.40167578384103586   0.6531927542415966   0.18344060507814625   0.38299025226421785   0.33959947485097086   0.15219273281664827   0.5275453226354317   0.32803973323074004   0.333194408851689   0.48687039293142514   0.41591158004222184   0.46314623887006867   0.3371287134262413   0.28509287148470325   0.018122035280359876   0.19484943089318074   0.8644877249214667   0.19133281862112506   0.9905768557446977   0.22036472411288013   0.8292835613344942   0.8600245286399116   0.0886609828842338   0.6568643731305565   0.42760777749345835   0.20683177439831507   0.9052203778060876   0.2738741208663386   0.08800830264248749   0.0546390415816668   0.3776750551706558   0.9458343876355986   0.7548138937907986   0.5677686486502417
0.961763475128434   0.4826881487655299   0.4176851803645572   0.2826757771655384   0.9436414398480741   0.28783871787234916   0.5531974554430905   0.09134295854441334   0.9530645841033764   0.06747399375946904   0.7239138941085963   0.2313184299045017   0.8644036012191426   0.4106096206289126   0.2963061166151379   0.024486655506186603   0.9591832234130551   0.136735499762574   0.2082978139726504   0.9698476139245198   0.5815081682423993   0.19090111212697541   0.4534839201818519   0.40207896527427817   0.6197446931139653   0.7082129633614455   0.03579873981729466   0.11940318810873977   0.6761032532658912   0.4203742454890963   0.4826012843742042   0.02806022956432644   0.7230386691625148   0.35290025172962725   0.7586873902656079   0.7967417996598247   0.8586350679433722   0.9422906311007146   0.46238127365047005   0.7722551441536382   0.8994518445303172   0.8055551313381407   0.25408345967781965   0.8024075302291184   0.317943676287918   0.6146540192111652   0.8005995394959677   0.4003285649548402   0.6981989831739527   0.9064410558497198   0.7648007996786731   0.2809253768461004   0.022095729908061534   0.48606681036062344   0.2821995153044689   0.25286514728177395   0.2990570607455467   0.1331665586309962   0.523512125038861   0.4561233476219492   0.44042199280217453   0.19087592753028154   0.06113085138839095   0.683868203468311
0.5409701482718573   0.3853207961921409   0.8070473917105713   0.8814606732391927   0.22302647198393935   0.7706667769809756   0.006447852214603546   0.48113210828435254   0.5248274888099866   0.8642257211312558   0.24164705253593044   0.20020673143825213   0.5027317589019251   0.37815891077063235   0.9594475372314616   0.9473415841564782   0.2036746981563784   0.24499235213963616   0.43593541219260057   0.49121823653452895   0.7632527053542039   0.054116424609354626   0.3748045608042096   0.8073500330662179   0.22228255708234657   0.6687956284172137   0.5677571690936383   0.9258893598270252   0.9992560850984072   0.8981288514362382   0.5613093168790347   0.44475725154267265   0.47442859628842055   0.03390313030498237   0.3196622643431043   0.24455052010442055   0.9716968373864954   0.65574421953435   0.36021472711164276   0.2972089359479424   0.768022139230117   0.41075186739471387   0.9242793149190422   0.8059906994134135   0.004769433875913118   0.35663544278535925   0.5494747541148326   0.9986406663471956   0.7824868767935665   0.6878398143681455   0.9817175850211943   0.07275130652017038   0.7832307916951594   0.7897109629319073   0.4204082681421596   0.6279940549774977   0.30880219540673887   0.755807832626925   0.1007460037990553   0.38344353487307714   0.33710535802024344   0.1000636130925749   0.7405312766874126   0.08623459892513473
0.5690832187901265   0.689311745697861   0.8162519617683703   0.2802438995117213   0.5643137849142134   0.3326763029125018   0.2667772076535377   0.2816032331645257   0.7818269081206468   0.6448364885443564   0.28505962263234336   0.2088519266443553   0.9985961164254874   0.855125525612449   0.8646513544901838   0.5808578716668577   0.6897939210187486   0.0993176929855241   0.7639053506911285   0.19741433679378048   0.3526885629985051   0.9992540798929492   0.023374074003715932   0.11117973786864575   0.7836053442083786   0.30994233419508815   0.2071221122353456   0.8309358383569245   0.21929155929416527   0.9772660312825864   0.9403449045818079   0.5493326051923988   0.4374646511735185   0.33242954273823005   0.6552852819494646   0.3404806785480435   0.43886853474803106   0.477304017125781   0.7906339274592807   0.7596228068811859   0.7490746137292825   0.3779863241402569   0.0267285767681523   0.5622084700874054   0.39638605073077743   0.3787322442473077   0.0033545027644363646   0.4510287322187596   0.6127807065223988   0.06878991005221954   0.7962323905290908   0.6200928938618351   0.3934891472282335   0.09152387876963318   0.8558874859472828   0.07076028866943632   0.9560244960547151   0.7590943360314032   0.2006022039978183   0.7302796101213929   0.517155961306684   0.2817903189056221   0.4099682765385375   0.9706568032402071
0.7680813475774014   0.9038039947653652   0.38323969977038524   0.4084483331528017   0.371695296846624   0.5250717505180575   0.37988519700594886   0.9574196009340421   0.7589145903242251   0.45628184046583803   0.5836528064768581   0.33732670707220697   0.3654254430959917   0.36475796169620484   0.7277653205295753   0.2665664184027707   0.4094009470412766   0.6056636256648017   0.527163116531757   0.5362868082813778   0.8922449857345927   0.3238733067591795   0.11719483999321943   0.5656300050411708   0.1241636381571912   0.4200693119938143   0.7339551402228341   0.15718167188836907   0.7524683413105672   0.8949975614757567   0.35406994321688534   0.19976207095432696   0.993553750986342   0.43871572100991874   0.7704171367400272   0.8624353638821199   0.6281283078903503   0.07395775931371393   0.042651816210451936   0.5958689454793493   0.21872736084907374   0.46829413364891226   0.5154886996786949   0.059582137197971514   0.3264823751144811   0.1444208268897327   0.39829385968547554   0.4939521321568007   0.2023187369572899   0.7243515148959184   0.6643387194626413   0.33677046026843166   0.44985039564672274   0.8293539534201617   0.31026877624575605   0.1370083893141047   0.4562966446603807   0.3906382324102429   0.5398516395057288   0.2745730254319847   0.8281683367700304   0.316680473096529   0.4971998232952769   0.6787040799526354
0.6094409759209567   0.8483863394476168   0.981711123616582   0.6191219427546639   0.28295860080647556   0.7039655125578841   0.5834172639311064   0.12516981059786314   0.08063986384918564   0.9796139976619657   0.919078544468465   0.7883993503294314   0.630789468202463   0.15026004424180395   0.6088097682227089   0.6513909610153268   0.17449282354208218   0.759621811831561   0.06895812871698016   0.3768179355833421   0.3463244867720518   0.442941338735032   0.5717583054217033   0.6981138556307067   0.7368835108510952   0.5945549992874153   0.5900471818051214   0.07899191287604279   0.4539249100446196   0.8905894867295312   0.0066299178740149714   0.9538221022781797   0.37328504619543396   0.9109754890675655   0.08755137340554996   0.1654227519487482   0.7424955779929711   0.7607154448257617   0.478741605182841   0.5140317909334214   0.5680027544508889   0.0010936329942006437   0.40978347646586083   0.13721385535007935   0.22167826767883705   0.5581522942591687   0.8380251710441575   0.4390999997193727   0.4847947568277419   0.9635972949717534   0.2479779892390362   0.3601080868433299   0.03086984678312233   0.0730078082422222   0.24134807136502123   0.40628598456515025   0.6575848005876884   0.1620323191746566   0.15379669795947126   0.24086323261640202   0.9150892225947174   0.40131687434889496   0.6750550927766303   0.7268314416829806
0.3470864681438285   0.40022324135469434   0.2652716163107695   0.5896175863329013   0.12540820046499146   0.8420709470955257   0.427246445266612   0.15051758661352857   0.6406134436372495   0.8784736521237723   0.17926845602757577   0.7904094997701987   0.6097435968541272   0.8054658438815501   0.9379203846625546   0.38412351520504845   0.9521587962664388   0.6434335247068934   0.7841236867030833   0.14326028258864643   0.037069573671721465   0.2421166503579985   0.10906859392645295   0.41642884090566584   0.689983105527893   0.8418934090033042   0.8437969776156834   0.8268112545727646   0.5645749050629015   0.9998224619077786   0.41655053234907147   0.676293667959236   0.9239614614256519   0.12134880978400625   0.23728207632149573   0.8858841681890374   0.3142178645715248   0.3158829659024562   0.2993616916589412   0.5017606529839889   0.36205906830508594   0.6724494411955627   0.5152380049558579   0.35850037039534244   0.3249894946333645   0.4303327908375642   0.40616941102940496   0.9420715294896767   0.6350063891054716   0.58843938183426   0.5623724334137216   0.11526027491691204   0.07043148404257002   0.5886169199264815   0.14582190106465004   0.43896660695767603   0.14647002261691805   0.46726811014247527   0.9085398247431543   0.5530824387686387   0.8322521580453933   0.15138514424001906   0.6091781330842131   0.051321785784649875
0.4701930897403073   0.4789357030444564   0.09394012812835519   0.6928214153893074   0.1452035951069428   0.04860291220689216   0.6877707170989502   0.7507498858996309   0.5101972060014712   0.46016353037263213   0.12539828368522868   0.6354896109827188   0.43976572195890123   0.8715466104461507   0.9795763826205787   0.19652300402504275   0.2932956993419832   0.4042785003036754   0.07103655787742431   0.643440565256404   0.4610435412965899   0.2528933560636563   0.4618584247932112   0.5921187794717542   0.9908504515562826   0.7739576530191999   0.367918296664856   0.8992973640824466   0.8456468564493398   0.7253547408123078   0.6801475795659058   0.14854747818281586   0.3354496504478685   0.26519121043967564   0.5547492958806771   0.513057867200097   0.8956839284889673   0.393644599993525   0.5751729132600985   0.3165348631750543   0.6023882291469841   0.9893660996898496   0.5041363553826742   0.6730942979186503   0.14134468785039414   0.7364727436261933   0.04227793058946299   0.08097551844689616   0.15049423629411152   0.9625150906069934   0.674359633924607   0.18167815436444948   0.3048473798447717   0.2371603497946855   0.9942120543587012   0.03313067618163361   0.9693977293969032   0.9719691393550098   0.4394627584780241   0.5200728089815365   0.07371380090793589   0.5783245393614848   0.8642898452179255   0.2035379458064822
0.4713255717609518   0.5889584396716352   0.36015348983525136   0.5304436478878319   0.3299808839105577   0.8524856960454419   0.3178755592457884   0.4494681294409358   0.17948664761644617   0.8899706054384486   0.6435159253211814   0.2677899750764863   0.8746392677716744   0.6528102556437632   0.6493038709624802   0.23465929889485268   0.9052415383747713   0.6808411162887533   0.20984111248445614   0.7145864899133162   0.8315277374668354   0.10251657692726848   0.34555126726653057   0.5110485441068339   0.3602021657058836   0.5135581372556333   0.9853977774312792   0.980604896219002   0.030221281795325898   0.6610724412101914   0.6675222181854908   0.5311367667780662   0.8507346341788797   0.7711018357717427   0.0240062928643094   0.26334679170157993   0.9760953664072053   0.11829158012797962   0.3747024219018292   0.028687492806727263   0.07085382803243401   0.4374504638392263   0.16486130941737304   0.31410100289341114   0.23932609056559861   0.33493388691195786   0.8193100421508425   0.8030524587865772   0.879123924859715   0.8213757496563245   0.8339122647195633   0.8224475625675752   0.8489026430643891   0.16030330844613322   0.16639004653407247   0.29131079578950897   0.9981680088855094   0.3892014726743905   0.14238375366976305   0.027964004087929026   0.022072642478304122   0.27090989254641085   0.7676813317679338   0.9992765112812018
0.9512188144458701   0.8334594287071845   0.6028200223505609   0.6851755083877906   0.7118927238802715   0.4985255417952266   0.7835099801997184   0.8821230496012135   0.8327687990205564   0.677149792138902   0.9495977154801551   0.059675487033638216   0.9838661559561673   0.5168464836927689   0.7832076689460826   0.7683646912441292   0.985698147070658   0.1276450110183784   0.6408239152763195   0.7404006871562002   0.9636255045923537   0.8567351184719676   0.8731425835083857   0.7411241758749985   0.012406690146483672   0.023275689764783076   0.2703225611578249   0.05594866748720782   0.3005139662662122   0.5247501479695564   0.48681258095810653   0.1738256178859944   0.4677451672456557   0.8476003558306543   0.5372148654779514   0.11415013085235617   0.48387901128948835   0.3307538721378855   0.7540071965318688   0.34578543960822694   0.49818086421883045   0.20310886111950707   0.11318328125554918   0.6053847524520267   0.5345553596264767   0.3463737426475395   0.24004069774716344   0.8642605765770283   0.5221486694799929   0.3230980528827564   0.9697181365893386   0.8083119090898204   0.22163470321378081   0.7983479049132   0.482905555631232   0.634486291203826   0.7538895359681251   0.9507475490825457   0.9456906901532806   0.5203361603514699   0.27001052467863673   0.6199936769446601   0.1916834936214118   0.17455072074324293
0.7718296604598063   0.4168848158251531   0.07850021236586262   0.5691659682912162   0.23727430083332965   0.0705110731776136   0.8384595146186992   0.704905391714188   0.7151256313533366   0.7474130202948572   0.8687413780293607   0.8965934826243676   0.4934909281395558   0.9490651153816572   0.38583582239812864   0.2621071914205415   0.7396013921714307   0.9983175662991115   0.4401451322448481   0.7417710310690717   0.46959086749279394   0.3783238893544514   0.24846163862343626   0.5672203103258288   0.6977612070329876   0.9614390735292982   0.16996142625757363   0.9980543420346125   0.460486906199658   0.8909280003516847   0.33150191163887444   0.29314895032042454   0.7453612748463213   0.1435149800568275   0.4627605336095138   0.396555467696057   0.2518703467067655   0.1944498646751703   0.07692471121138518   0.13444827627551548   0.5122689545353348   0.19613229837605878   0.6367795789665371   0.3926772452064438   0.0426780870425409   0.8178084090216073   0.38831794034310085   0.8254569348806151   0.3449168800095533   0.8563693354923091   0.21835651408552723   0.8274025928460025   0.8844299738098953   0.9654413351406244   0.8868546024466527   0.5342536425255779   0.13906869896357396   0.8219263550837969   0.42409406883713896   0.137698174829521   0.8871983522568084   0.6274764904086266   0.34716935762575374   0.003249898554005523
0.3749293977214736   0.4313441920325678   0.7103897786592166   0.6105726533475617   0.3322513106789327   0.6135357830109605   0.3220718383161158   0.7851157184669466   0.9873344306693794   0.7571664475186514   0.10371532423058857   0.9577131256209441   0.10290445685948414   0.7917251123780269   0.2168607217839358   0.42345948309536613   0.9638357578959103   0.96979875729423   0.7927666529467968   0.28576130826584517   0.07663740563910176   0.34232226688560347   0.4455972953210431   0.28251140971183963   0.7017080079176281   0.9109780748530356   0.7352075166618265   0.6719387563642779   0.36945669723869545   0.2974422918420752   0.4131356783457107   0.8868230378973312   0.382122266569316   0.5402758443234239   0.3094203541151221   0.9291099122763871   0.2792178097098319   0.7485507319453969   0.09255963233118629   0.505650429181021   0.3153820518139217   0.7787519746511669   0.2997929793843894   0.21988912091517582   0.2387446461748199   0.4364297077655634   0.8541956840633463   0.9373777112033362   0.5370366382571917   0.5254516329125277   0.11898816740151985   0.2654389548390583   0.1675799410184963   0.22800934107045254   0.7058524890558092   0.3786159169417271   0.7854576744491802   0.6877334967470287   0.3964321349406871   0.44950600466533996   0.5062398647393485   0.9391827648016318   0.30387250260950077   0.943855575484319
0.19085781292542672   0.1604307901504649   0.004079523225111354   0.7239664545691432   0.9521131667506069   0.7240010823849015   0.14988383916176504   0.786588743365807   0.41507652849341503   0.19854944947237377   0.030895671760245186   0.5211497885267486   0.24749658747491876   0.9705401084019212   0.325043182704436   0.1425338715850216   0.46203891302573846   0.2828066116548925   0.9286110477637489   0.6930278669196817   0.9557990482863901   0.34362384685326075   0.6247385451542482   0.7491722914353627   0.7649412353609634   0.18319305670279587   0.6206590219291368   0.025205836866219487   0.8128280686103565   0.4591919743178944   0.4707751827673718   0.23861709350041252   0.39775154011694147   0.2606425248455206   0.4398795110071266   0.7174673049736638   0.1502549526420227   0.2901024164435994   0.11483632830269057   0.5749334333886422   0.6882160396162842   0.0072958047887068484   0.18622528053894163   0.8819055664689607   0.7324169913298941   0.6636719579354461   0.5614867353846935   0.13273327503359797   0.9674757559689309   0.48047890123265025   0.9408277134555567   0.10752743816737849   0.15464768735857434   0.021286926914755866   0.4700525306881849   0.8689103446669659   0.7568961472416329   0.7606444020692352   0.030173019681058334   0.15144303969330208   0.6066411945996102   0.4705419856256359   0.9153366913783677   0.5765096063046599
0.9184251549833259   0.46324618083692903   0.7291114108394261   0.6946040398356992   0.18600816365343176   0.799574222901483   0.16762467545473264   0.5618707648021012   0.2185324076845009   0.31909532166883275   0.22679696199917596   0.4543433266347227   0.06388472032592657   0.2978083947540769   0.756744431310991   0.5854329819677567   0.3069885730842937   0.5371639926848416   0.7265714116299327   0.4339899422744547   0.7003473784846835   0.0666220070592057   0.811234720251565   0.8574803359697949   0.7819222235013576   0.6033758262222767   0.08212330941213883   0.16287629613409565   0.5959140598479259   0.8038016033207938   0.9144986339574062   0.6010055313319944   0.37738165216342495   0.484706281651961   0.6877016719582302   0.1466622046972717   0.3134969318374984   0.1868978868978841   0.9309572406472392   0.5612292227295149   0.006508358753204675   0.6497338942130425   0.20438582901730645   0.12723928045506025   0.3061609802685211   0.5831118871538368   0.3931511087657415   0.2697589444852654   0.5242387567671636   0.9797360609315602   0.3110277993536027   0.10688264835116974   0.9283246969192377   0.1759344576107664   0.3965291653961965   0.5058771170191753   0.5509430447558127   0.6912281759588054   0.7088274934379662   0.3592149123219036   0.23744611291831436   0.5043302890609213   0.7778702527907271   0.7979856895923887
0.23093775416510967   0.8545963948478787   0.5734844237734206   0.6707464091373284   0.9247767738965885   0.271484507694042   0.1803333150076791   0.40098746465206303   0.400538017129425   0.2917484467624818   0.8693055156540764   0.2941048163008933   0.4722133202101873   0.11581398915171541   0.47277635025787995   0.788227699281718   0.9212702754543746   0.42458581319291   0.7639488568199138   0.4290127869598144   0.6838241625360603   0.9202555241319887   0.9860786040291867   0.6310270973674257   0.45288640837095057   0.06565912928410993   0.41259418025576605   0.9602806882300973   0.528109634474362   0.794174621590068   0.23226086524808695   0.5592932235780342   0.12757161734493702   0.5024261748275861   0.36295534959401055   0.26518840727714094   0.6553582971347497   0.38661218567587075   0.8901789993361305   0.47696070799542295   0.7340880216803751   0.9620263724829607   0.12623014251621686   0.047947921035608534   0.050263859144314874   0.04177084835097208   0.14015153848703021   0.41692082366818284   0.5973774507733643   0.9761117190668621   0.7275573582312642   0.45664013543808557   0.06926781629900226   0.18193709747679418   0.49529649298317724   0.8973469118600513   0.9416961989540652   0.679510922649208   0.13234114338916672   0.6321585045829103   0.2863379018193155   0.2928987369733373   0.24216214405303615   0.15519779658748747
0.5522498801389404   0.3308723644903765   0.11593200153681928   0.10724987555187893   0.5019860209946255   0.28910151613940444   0.975780463049789   0.6903290518836961   0.9046085702212613   0.31298979707254226   0.2482231048185249   0.23368891644561054   0.8353407539222589   0.1310526995957481   0.7529266118353476   0.33634200458555924   0.8936445549681937   0.4515417769465401   0.6205854684461809   0.7041835000026488   0.6073066531488782   0.1586430399732028   0.37842332439314474   0.5489857034151614   0.05505677300993779   0.8277706754828263   0.2624913228563255   0.44173582786328247   0.5530707520153122   0.5386691593434219   0.28671085980653643   0.7514067759795864   0.648462181794051   0.2256793622708796   0.038487754988011554   0.5177178595339758   0.8131214278717921   0.09462666267513148   0.2855611431526639   0.18137585494841654   0.9194768729035983   0.6430848857285915   0.664975674706483   0.4771923549457677   0.3121702197547201   0.4844418457553886   0.28655235031333826   0.9282066515306063   0.2571134467447823   0.6566711702725623   0.024061027457012746   0.4864708236673239   0.7040426947294701   0.11800201092914042   0.7373501676504763   0.7350640476877376   0.05558051293541906   0.8923226486582608   0.6988624126624647   0.21734618815376178   0.242459085063627   0.7976959859831293   0.41330126950980084   0.03597033320534522
0.3229822121600287   0.15461110025453795   0.7483255948033178   0.5587779782595775   0.01081199240530861   0.6701692544991493   0.46177324448997964   0.6305713267289712   0.7536985456605263   0.013498084226587055   0.43771221703296687   0.1441005030616473   0.049655850931056233   0.8954960732974466   0.7003620493824906   0.40903645537390976   0.9940753379956372   0.0031734246391857935   0.0014996367200257837   0.19169026722014798   0.7516162529320102   0.20547743865605644   0.5881983672102249   0.15571993401480275   0.4286340407719814   0.050866338401518496   0.839872772406907   0.5969419557552252   0.41782204836667286   0.38069708390236917   0.37809952791692747   0.966370629026254   0.6641235027061465   0.36719899967578207   0.9403873108839605   0.8222701259646068   0.6144676517750903   0.47170292637833544   0.24002526150147002   0.41323367059069704   0.6203923137794531   0.46852950173914965   0.23852562478144423   0.22154340337054906   0.868776060847443   0.2630520630830932   0.6503272575712193   0.0658234693557463   0.4401420200754615   0.21218572468157473   0.8104544851643123   0.46888151360052105   0.02231997170878869   0.8314886407792056   0.43235495724738476   0.502510884574267   0.3581964690026421   0.46428964110342347   0.4919676463634242   0.6802407586096602   0.7437288172275519   0.9925867147250881   0.2519423848619542   0.26700708801896317
0.12333650344809872   0.5240572129859383   0.01341676008050993   0.04546368464841412   0.25456044260065575   0.2610051499028451   0.3630895025092906   0.9796402152926679   0.8144184225251943   0.048819425221270404   0.5526350173449783   0.5107587016921468   0.7920984508164055   0.21733078444206483   0.1202800600975936   0.00824781711787978   0.4339019818137634   0.7530411433386414   0.6283124137341694   0.3280070585082196   0.6901731645862116   0.7604544286135533   0.3763700288722152   0.0609999704892564   0.5668366611381128   0.23639721562761495   0.3629532687917053   0.015536285840842287   0.3122762185374571   0.9753920657247698   0.9998637662824147   0.03589607054817447   0.4978577960122628   0.9265726405034994   0.4472287489374363   0.5251373688560277   0.7057593451958573   0.7092418560614346   0.3269486888398427   0.5168895517381479   0.2718573633820938   0.9562007127227933   0.6986362751056733   0.18888249322992834   0.5816841987958823   0.19574628410923994   0.32226624623345806   0.12788252274067194   0.014847537657769475   0.959349068481625   0.9593129774417528   0.11234623689982966   0.7025713191203125   0.9839570027568552   0.9594492111593381   0.07645016635165519   0.2047135231080496   0.05738436225335579   0.5122204622219018   0.5513127974956274   0.4989541779121924   0.3481425061919212   0.1852717733820591   0.03442324575747956
0.22709681453009853   0.39194179346912794   0.4866354982763858   0.8455407525275512   0.6454126157342163   0.196195509359888   0.16436925204292774   0.7176582297868792   0.6305650780764468   0.23684644087826298   0.20505627460117495   0.6053119928870496   0.9279937589561343   0.2528894381214078   0.24560706344183686   0.5288618265353944   0.7232802358480848   0.195505075868052   0.733386601219935   0.9775490290397669   0.22432605793589236   0.8473625696761308   0.5481148278378759   0.9431257832822874   0.9972292434057938   0.45542077620700283   0.061479329561490124   0.09758503075473614   0.3518166276715776   0.25922526684711483   0.8971100775185624   0.37992680096785686   0.7212515495951308   0.02237882596885188   0.6920538029173874   0.7746148080808073   0.7932577906389965   0.7694893878474441   0.4464467394755506   0.2457529815454129   0.0699775547909118   0.5739843119793921   0.7130601382556155   0.268203952505646   0.8456514968550195   0.7266217423032613   0.1649453104177396   0.32507816922335864   0.8484222534492256   0.2712009660962585   0.10346598085624947   0.22749313846862249   0.49660562577764805   0.01197569924914361   0.20635590333768708   0.8475663375007656   0.7753540761825172   0.9895968732802918   0.5143021004202997   0.0729515294199583   0.9820962855435207   0.22010748543284764   0.06785536094474907   0.8271985478745454
0.9121187307526089   0.6461231734534555   0.35479522268913355   0.5589945953688995   0.0664672338975894   0.9195014311501942   0.18984991227139394   0.23391642614554084   0.2180449804483638   0.6483004650539358   0.08638393141514446   0.0064232876769183605   0.7214393546707157   0.6363247658047921   0.8800280280774574   0.15885695017615278   0.9460852784881986   0.6467278925245004   0.3657259276571577   0.08590542075619446   0.9639889929446779   0.4266204070916528   0.29787056671240864   0.25870687288164906   0.05187026219206902   0.7804972336381972   0.9430753440232751   0.6997122775127496   0.9854030282944796   0.860995802488003   0.7532254317518812   0.46579585136720875   0.7673580478461158   0.2126953374340673   0.6668415003367367   0.4593725636902904   0.045918693175400094   0.5763705716292752   0.7868134722592793   0.30051561351413764   0.09983341468720154   0.9296426791047747   0.4210875446021216   0.21461019275794316   0.13584442174252365   0.503022272013122   0.123216977889713   0.9559033198762941   0.08397415955045463   0.7225250383749248   0.18014163386643792   0.2561910423635445   0.09857113125597503   0.8615292358869218   0.4269162021145568   0.7903951909963357   0.33121308340985917   0.6488338984528544   0.7600747017778201   0.33102262730604537   0.28529439023445907   0.07246332682357927   0.9732612295185407   0.030507013791907723
0.18546097554725757   0.1428206477188045   0.552173684916419   0.8158968210339645   0.04961655380473391   0.6397983757056825   0.4289567070267061   0.8599935011576705   0.9656423942542792   0.9172733373307578   0.24881507316026816   0.603802458794126   0.8670712629983043   0.055744101443836076   0.8218988710457114   0.8134072677977902   0.5358581795884451   0.40691020299098163   0.061824169267891346   0.4823846404917448   0.250563789353986   0.3344468761674024   0.08856293974935063   0.4518776266998371   0.0651028138067284   0.19162622844859786   0.5363892548329315   0.6359808056658726   0.015486260001994493   0.5518278527429153   0.10743254780622548   0.7759873045082021   0.04984386574771522   0.6345545154121576   0.8586174746459573   0.17218484571407616   0.18277260274941096   0.5788104139683214   0.03671860360024591   0.358777577916286   0.6469144231609659   0.17190021097733982   0.9748944343323546   0.8763929374245412   0.39635063380697994   0.8374533348099374   0.886331494583004   0.4245153107247041   0.33124782000025155   0.6458271063613396   0.3499422397500724   0.7885345050588316   0.31576155999825706   0.09399925361842427   0.2425096919438469   0.012547200550629509   0.2659176942505418   0.45944473820626675   0.3838922172978896   0.8403623548365533   0.08314509150113085   0.8806343242379453   0.34717361369764366   0.48158477692026735
0.43623066834016494   0.7087341132606054   0.3722791793652891   0.6051918394957261   0.03988003453318503   0.8712807784506681   0.48594768478228517   0.18067652877102203   0.7086322145329335   0.22545367208932846   0.1360054450322128   0.3921420237121904   0.39287065453467646   0.13145441847090417   0.8934957530883659   0.3795948231615609   0.12695296028413466   0.6720096802646375   0.5096035357904763   0.5392324683250076   0.043807868783003794   0.7913753560266922   0.16242992209283266   0.057647691404740235   0.6075772004428388   0.08264124276608667   0.7901507427275436   0.4524558519090141   0.5676971659096538   0.21136046431541863   0.30420305794525837   0.2717793231379921   0.8590649513767203   0.9859067922260901   0.1681976129130456   0.8796372994258017   0.46619429684204383   0.854452373755186   0.2747018598246797   0.5000424762642407   0.33924133655790917   0.18244269349054856   0.7650983240342034   0.9608100079392332   0.29543346777490537   0.3910673374638564   0.6026684019413707   0.903162316534493   0.6878562673320665   0.30842609469776977   0.8125176592138271   0.45070646462547886   0.12015910142241275   0.09706563038235112   0.5083146012685688   0.17892714148748676   0.2610941500456924   0.11115883815626094   0.3401169883555232   0.29928984206168513   0.7948998532036486   0.2567064644010749   0.06541512853084347   0.7992473657974444
0.4556585166457394   0.07426377091052638   0.30031680449664006   0.8384373578582112   0.16022504887083405   0.68319643344667   0.6976484025552694   0.9352750413237182   0.4723687815387675   0.3747703387489002   0.8851307433414421   0.4845685766982394   0.35220968011635473   0.2777047083665491   0.37681614207287345   0.3056414352107526   0.09111553007066231   0.16654587021028816   0.036699153717350254   0.006351593149067513   0.2962156768670137   0.9098394058092132   0.9712840251865068   0.20710422735162315   0.8405571602212742   0.8355756348986868   0.6709672206898667   0.368666869493412   0.6803321113504402   0.15237920145201686   0.9733188181345973   0.43339182816969374   0.20796332981167276   0.7776088627031167   0.08818807479315516   0.9488232514714544   0.855753649695318   0.49990415433656754   0.7113719327202818   0.6431818162607017   0.7646381196246557   0.3333582841262794   0.6746727790029314   0.6368302231116343   0.468422442757642   0.42351887831706614   0.7033887538164247   0.4297259957600111   0.6278652825363678   0.5879432434183793   0.03242153312655798   0.0610591262665991   0.9475331711859275   0.43556404196636245   0.059102714991960625   0.6276672980969054   0.7395698413742547   0.6579551792632459   0.9709146401988055   0.678844046625451   0.8838161916789368   0.1580510249266783   0.2595427074785237   0.03566223036474923
0.11917807205428103   0.8246927408003989   0.5848699284755923   0.39883200725311496   0.650755629296639   0.40117386248333275   0.8814811746591675   0.9691060114931039   0.022890346760271338   0.8132306190649534   0.8490596415326096   0.9080468852265048   0.07535717557434388   0.37766657709859097   0.789956926540649   0.28037958712959943   0.33578733420008916   0.7197113978353452   0.8190422863418435   0.6015355405041485   0.45197114252115245   0.5616603729086669   0.5594995788633198   0.5658733101393992   0.3327930704668714   0.736967632108268   0.9746296503877275   0.16704130288628424   0.6820374411702324   0.3357937696249352   0.09314847572855994   0.19793529139318036   0.659147094409961   0.5225631505599817   0.24408883419595037   0.28988840616667555   0.5837899188356171   0.1448965734613907   0.4541319076553014   0.009508819037076094   0.248002584635528   0.4251851756260455   0.6350896213134579   0.40797327853292764   0.7960314421143756   0.8635248027173786   0.07559004245013816   0.8420999683935284   0.46323837164750414   0.1265571706091107   0.10096039206241066   0.6750586655072441   0.7812009304772718   0.7907634009841755   0.007811916333850706   0.47712337411406375   0.12205383606731075   0.2682002504241938   0.7637230821379003   0.18723496794738823   0.5382639172316936   0.12330367696280312   0.30959117448259893   0.17772614891031213
0.2902613325961656   0.6981185013367576   0.674501553169141   0.7697528703773845   0.49422989048179006   0.8345936986193789   0.5989115107190028   0.9276529019838561   0.03099151883428588   0.7080365280102682   0.4979511186565922   0.252594236476612   0.2497905883570141   0.9172731270260926   0.4901392023227415   0.7754708623625483   0.12773675228970335   0.6490728766018988   0.7264161201848411   0.58823589441516   0.5894728350580097   0.5257691996390957   0.4168249457022422   0.41050974550484787   0.29921150246184414   0.8276506983023382   0.7423233925331012   0.6407568751274634   0.8049816119800541   0.9930569996829592   0.14341188181409836   0.7131039731436073   0.7739900931457683   0.285020471672691   0.6454607631575062   0.46050973666699524   0.5241995047887541   0.36774734464659836   0.15532156083476473   0.685038874304447   0.39646275249905083   0.7186744680446995   0.4289054406499236   0.09680297988928699   0.8069899174410411   0.1929052684056038   0.012080494947681384   0.6862932343844391   0.5077784149791968   0.3652545701032656   0.2697571024145802   0.04553635925697573   0.7027968029991427   0.3721975704203064   0.12634522060048178   0.3324323861133685   0.9288067098533745   0.08717709874761535   0.4808844574429756   0.8719226494463732   0.40460720506462033   0.719429754101017   0.32556289660821086   0.18688377514192625
0.008144452565569539   0.000755286056317455   0.8966574559582873   0.09008079525263928   0.2011545351245285   0.8078500176507136   0.8845769610106059   0.40378756086820017   0.6933761201453316   0.44259544754744806   0.6148198585960257   0.3582512016112244   0.9905793171461889   0.07039787712714166   0.4884746379955439   0.025818815497855956   0.06177260729281434   0.9832207783795263   0.007590180552568329   0.1538961660514827   0.657165402228194   0.2637910242785093   0.6820272839443574   0.9670123909095565   0.6490209496626245   0.2630357382221919   0.7853698279860701   0.8769315956569171   0.44786641453809595   0.4551857205714782   0.9007928669754643   0.47314403478871697   0.7544902943927644   0.01259027302403017   0.28597300837943856   0.11489283317749253   0.7639109772465755   0.9421923958968885   0.7974983703838946   0.08907401767963657   0.7021383699537612   0.9589716175173623   0.7899081898313263   0.9351778516281539   0.044972967725567185   0.6951805932388528   0.10788090588696886   0.9681654607185974   0.3959520180629427   0.432144855016661   0.32251107790089867   0.0912338650616803   0.9480856035248467   0.9769591344451828   0.4217182109254344   0.6180898302729633   0.1935953091320824   0.9643688614211526   0.1357452025459958   0.5031969970954707   0.42968433188550686   0.022176465524264128   0.33824683216210116   0.4141229794158342
0.7275459619317457   0.06320484800690192   0.5483386423307749   0.47894512778768034   0.6825729942061785   0.368024254768049   0.440457736443806   0.5107796670690828   0.2866209761432358   0.935879399751388   0.11794665854290731   0.41954580200740255   0.338535372618389   0.9589202653062052   0.6962284476174729   0.8014559717344393   0.14494006348630664   0.9945514038850525   0.5604832450714772   0.2982589746389685   0.7152557316007998   0.9723749383607884   0.22223641290937596   0.8841359952231342   0.9877097696690541   0.9091700903538865   0.6738977705786011   0.40519086743545396   0.3051367754628756   0.5411458355858375   0.2334400341347951   0.8944112003663711   0.018515799319639856   0.6052664358344495   0.1154933755918878   0.4748653983589685   0.6799804267012508   0.6463461705282443   0.4192649279744149   0.6734094266245293   0.5350403632149442   0.6517947666431918   0.8587816829029378   0.3751504519855608   0.8197846316141444   0.6794198282824033   0.6365452699935618   0.4910144567624265   0.8320748619450904   0.7702497379285169   0.9626474994149606   0.08582358932697254   0.5269380864822147   0.2291039023426794   0.7292074652801656   0.19141238896060142   0.5084222871625749   0.6238374665082299   0.6137140896882778   0.7165469906016328   0.8284418604613241   0.9774912959799856   0.19444916171386287   0.04313756397710361
0.2934014972463798   0.3256965293367939   0.3356674788109251   0.6679871119915428   0.4736168656322354   0.6462767010543905   0.6991222088173633   0.1769726552291163   0.641542003687145   0.8760269631258737   0.7364747094024027   0.09114906590214376   0.1146039172049303   0.6469230607831943   0.0072672441222371605   0.8997366769415424   0.6061816300423555   0.023085594274964333   0.39355315443395944   0.18318968633990945   0.7777397695810314   0.04559429829497869   0.19910399272009655   0.14005212236280584   0.4843382723346516   0.7198977689581848   0.8634365139091714   0.472065010371263   0.010721406702416246   0.07362106790379427   0.16431430509180805   0.2950923551421467   0.36917940301527125   0.1975941047779206   0.4278395956894054   0.20394328924000296   0.25457548581034095   0.5506710439947263   0.4205723515671682   0.30420661229846063   0.6483938557679855   0.5275854497197621   0.027019197133208776   0.12101692595855118   0.8706540861869541   0.4819911514247833   0.8279152044131122   0.9809648035957453   0.38631581385230246   0.7620933824665985   0.9644786905039407   0.5088997932244823   0.37559440714988623   0.6884723145628042   0.8001643854121328   0.2138074380823356   0.006415004134615012   0.4908782097848836   0.37232478972272737   0.009864148842332634   0.7518395183242741   0.9402071657901573   0.9517524381555592   0.705657536543872
0.10344566255628858   0.4126217160703953   0.9247332410223504   0.5846406105853208   0.23279157636933448   0.9306305646456119   0.09681803660923818   0.6036758069895755   0.846475762517032   0.1685371821790134   0.13233934610529738   0.09477601376509318   0.47088135536714576   0.48006486761620915   0.33217496069316466   0.8809685756827575   0.46446635123253077   0.9891866578313255   0.9598501709704372   0.871104426840425   0.7126268329082567   0.04897949204116826   0.008097732814878071   0.16544689029655293   0.6091811703519681   0.636357775970773   0.08336449179252767   0.5808062797112321   0.3763895939826336   0.705727211325161   0.9865464551832894   0.9771304727216567   0.5299138314656016   0.5371900291461477   0.8542071090779921   0.8823544589565634   0.05903247609845583   0.057125161529938503   0.5220321483848275   0.001385883273805838   0.5945661248659251   0.06793850369861296   0.5621819774143902   0.13028145643338088   0.8819392919576684   0.0189590116574447   0.5540842445995121   0.9648345661368279   0.2727581216057003   0.3826012356866717   0.47071975280698447   0.38402828642559583   0.8963685276230667   0.6768740243615107   0.484173297623695   0.40689781370393924   0.3664546961574651   0.13968399521536295   0.6299661885457029   0.5245433547473758   0.30742222005900927   0.08255883368542447   0.10793404016087543   0.52315747147357
0.7128560951930842   0.014620329986811495   0.5457520627464852   0.3928760150401891   0.8309168032354158   0.9956613183293668   0.9916678181469731   0.42804144890336115   0.5581586816297155   0.6130600826426951   0.5209480653399886   0.0440131624777653   0.6617901540066488   0.9361860582811845   0.03677476771629365   0.637115348773826   0.2953354578491837   0.7965020630658215   0.40680857917059077   0.11257199402645028   0.9879132377901744   0.713943229380397   0.29887453900971533   0.5894145225528803   0.2750571425970902   0.6993228993935856   0.75312247626323   0.19653850751269125   0.4441403393616744   0.7036615810642187   0.761454658116257   0.7684970586093302   0.8859816577319589   0.09060149842152367   0.24050659277626832   0.7244838961315648   0.22419150372531008   0.1544154401403392   0.20373182505997467   0.08736854735773873   0.9288560458761264   0.3579133770745177   0.7969232458893839   0.9747965533312885   0.940942808085952   0.6439701476941206   0.4980487068796686   0.3853820307784081   0.6658856654888617   0.944647248300535   0.7449262306164385   0.18884352326571688   0.22174532612718736   0.24098566723631631   0.9834715725001816   0.42034646465638675   0.3357636683952285   0.15038416881479263   0.7429649797239133   0.695862568524822   0.11157216466991841   0.9959687286744534   0.5392331546639385   0.6084940211670832
0.18271611879379204   0.6380553515999358   0.7423099087745546   0.6336974678357948   0.24177331070784008   0.9940852039058151   0.244261201894886   0.24831543705738665   0.5758876452189784   0.04943795560528006   0.4993349712784475   0.05947191379166977   0.354142319091791   0.8084522883689638   0.5158633987782659   0.639125449135283   0.018378650696562526   0.6580681195541711   0.7728984190543526   0.943262880610461   0.9068064860266442   0.6620993908797177   0.23366526439041413   0.3347688594433778   0.724090367232852   0.024044039279781902   0.4913553556158595   0.701071391607583   0.482317056525012   0.02995883537396677   0.2470941537209735   0.45275595455019635   0.9064294113060336   0.9805208797686867   0.747759182442526   0.3932840407585266   0.5522870922142427   0.17206859139972297   0.23189578366426009   0.7541585916232436   0.5339084415176801   0.5140004718455519   0.4589973646099074   0.8108957110127826   0.627101955491036   0.8519010809658342   0.22533210021949326   0.47612685156940476   0.903011588258184   0.8278570416860523   0.7339767446036337   0.7750554599618217   0.4206945317331719   0.7978982063120855   0.4868825908826603   0.32229950541162533   0.5142651204271383   0.8173773265433988   0.7391234084401342   0.9290154646530987   0.9619780282128957   0.6453087351436758   0.5072276247758741   0.17485687302985514
0.4280695866952156   0.13130826329812398   0.048230260165966786   0.36396116201707257   0.8009676312041796   0.2794071823322898   0.8228981599464735   0.8878343104476678   0.8979560429459957   0.4515501406462375   0.08892141534283977   0.11277885048584611   0.4772615112128238   0.653651934334152   0.6020388244601795   0.7904793450742208   0.9629963907856856   0.8362746077907531   0.8629154160200453   0.861463880421122   0.0010183625727898235   0.19096587264707734   0.35568779124417105   0.6866070073912669   0.5729487758775742   0.059657609348953346   0.3074575310782043   0.3226458453741943   0.7719811446733946   0.7802504270166636   0.48455937113173075   0.4348115349265264   0.8740251017273989   0.32870028637042603   0.395637955788891   0.3220326844406803   0.3967635905145751   0.6750483520362741   0.7935991313287115   0.5315533393664595   0.4337671997288896   0.8387737442455209   0.9306837153086662   0.6700894589453376   0.43274883715609974   0.6478078715984436   0.5749959240644952   0.9834824515540707   0.8598000612785255   0.5881502622494902   0.2675383929862909   0.6608366061798764   0.08781891660513091   0.8078998352328267   0.7829790218545601   0.22602507125334997   0.21379381487773202   0.4791995488624006   0.38734106606566915   0.9039923868126697   0.817030224363157   0.8041511968261266   0.5937419347369577   0.37243904744621015
0.3832630246342673   0.9653774525806056   0.6630582194282915   0.7023495885008726   0.9505141874781676   0.31756958098216204   0.08806229536379624   0.7188671369468019   0.09071412619964205   0.7294193187326719   0.8205239023775054   0.05803053076692555   0.002895209594511128   0.9215194834998451   0.03754488052294524   0.8320054595135755   0.7891013947167791   0.44231993463744457   0.6502038144572762   0.9280130727009059   0.9720711703536222   0.638168737811318   0.056461879720318464   0.5555740252546958   0.5888081457193548   0.6727912852307124   0.39340366029202706   0.8532244367538231   0.6382939582411873   0.3552217042485503   0.30534136492823083   0.13435729980702116   0.5475798320415453   0.6258023855158785   0.48481746255072544   0.07632676904009562   0.5446846224470341   0.7042829020160334   0.4472725820277802   0.24432130952652006   0.755583227730255   0.2619629673785888   0.797068767570504   0.31630823682561415   0.7835120573766328   0.6237942295672708   0.7406068878501856   0.7607342115709185   0.19470391165727796   0.9510029443365584   0.3472032275581586   0.9075097748170953   0.5564099534160907   0.595781240088008   0.04186186262992777   0.7731524750100741   0.008830121374545493   0.9699788545721295   0.5570444000792023   0.6968257059699785   0.4641454989275114   0.2656959525560962   0.10977181805142211   0.45250439644345847
0.7085622711972565   0.003732985177507353   0.312703050480918   0.1361961596178443   0.9250502138206236   0.37993875561023654   0.5720961626307324   0.37546194804692584   0.7303463021633456   0.42893581127367814   0.2248929350725738   0.46795217322983057   0.17393634874725494   0.83315457118567   0.18303107244264602   0.6947996982197564   0.16510622737270944   0.8631757166135405   0.6259866723634437   0.9979739922497779   0.7009607284451981   0.5974797640574443   0.5162148543120216   0.5454695958063195   0.9923984572479416   0.593746778879937   0.2035118038311036   0.40927343618847517   0.067348243427318   0.21380802326970044   0.6314156412003712   0.03381148814154933   0.33700194126397237   0.7848722119960223   0.4065227061277974   0.5658593149117188   0.1630655925167174   0.9517176408103523   0.22349163368515138   0.8710596166919623   0.997959365144008   0.08854192419681173   0.5975049613217077   0.8730856244421844   0.29699863669880994   0.4910621601393674   0.08129010700968606   0.3276160286358649   0.3046001794508683   0.8973153812594304   0.8777783031785825   0.9183425924473897   0.2372519360235503   0.68350735798973   0.24636266197821124   0.8845311043058404   0.900249994759578   0.8986351459937076   0.8398399558504138   0.3186717893941216   0.7371844022428605   0.9469175051833554   0.6163483221652625   0.4476121727021593
0.7392250370988526   0.8583755809865437   0.01884336084355477   0.574526548259975   0.4422264004000427   0.3673134208471763   0.9375532538338687   0.24691051962411   0.1376262209491744   0.4699980395877459   0.05977495065528624   0.3285679271767203   0.9003742849256241   0.7864906815980159   0.813412288677075   0.4440368228708799   0.00012429016604613733   0.8878555356043083   0.9735723328266611   0.12536503347675831   0.26293988792318557   0.9409380304209528   0.35722401066139875   0.6777528607745991   0.523714850824333   0.08256244943440917   0.33838064981784394   0.10322631251462411   0.0814884504242903   0.7152490285872329   0.40082739598397527   0.8563157928905141   0.9438622294751159   0.245250988999487   0.341052445328689   0.5277478657137938   0.04348794454949182   0.4587603074014711   0.527640156651614   0.08371104284291389   0.04336365438344568   0.5709047717971628   0.5540678238249529   0.9583460093661555   0.7804237664602601   0.62996674137621   0.19684381316355412   0.2805931485915566   0.2567089156359271   0.5474042919418008   0.8584631633457102   0.17736683607693246   0.1752204652116368   0.8321552633545679   0.4576357673617349   0.32105104318641836   0.2313582357365209   0.5869042743550809   0.1165833220330459   0.7933031774726246   0.18787029118702908   0.1281439669536098   0.5889431653814319   0.7095921346297106
0.1445066368035834   0.5572391951564469   0.03487534155647904   0.751246125263555   0.3640828703433233   0.927272453780237   0.8380315283929249   0.47065297667199846   0.10737395470739619   0.3798681618384362   0.9795683650472148   0.293286140595066   0.9321534894957594   0.5477128984838683   0.5219325976854798   0.9722350974086477   0.7007952537592385   0.9608086241287874   0.40534927565243395   0.17893191993602314   0.5129249625722094   0.8326646571751776   0.8164061102710021   0.46933978530631254   0.368418325768626   0.2754254620187306   0.781530768714523   0.7180936600427574   0.0043354554253027065   0.3481530082384936   0.943499240321598   0.247440683370759   0.8969615007179065   0.9682848464000574   0.9639308752743834   0.954154542775693   0.9648080112221471   0.4205719479161891   0.4419982775889035   0.9819194453670453   0.26401275746290864   0.4597633237874017   0.03664900193646954   0.8029875254310221   0.7510877948906992   0.6270986666122241   0.22024289166546748   0.33364774012470966   0.3826694691220732   0.35167320459349355   0.43871212295094447   0.6155540800819521   0.3783340136967705   0.003520196354999967   0.49521288262934643   0.3681133967111932   0.48137251297886396   0.03523534995494258   0.5312820073549631   0.4139588539355002   0.5165645017567169   0.6146634020387535   0.0892837297660596   0.4320394085684549
0.2525517442938082   0.15490007825135177   0.05263472782959006   0.6290518831374328   0.501463949403109   0.5278014116391276   0.8323918361641226   0.2954041430127231   0.11879448028103581   0.17612820704563406   0.3936797132131781   0.679850062930771   0.7404604665842653   0.17260801069063408   0.8984668305838317   0.31173666621957774   0.2590879536054013   0.13737266073569152   0.3671848232288686   0.8977778122840776   0.7425234518486845   0.5227092586969381   0.277901093462809   0.46573840371562264   0.48997170755487623   0.36780918044558625   0.22526636563321895   0.8366865205781899   0.9885077581517672   0.8400077688064587   0.39287452946909635   0.5412823775654668   0.8697132778707314   0.6638795617608246   0.9991948162559183   0.8614323146346958   0.12925281128646607   0.4912715510701905   0.10072798567208661   0.5496956484151181   0.8701648576810648   0.35389889033449895   0.733543162443218   0.6519178361310405   0.12764140583238026   0.831189631637561   0.455642068980409   0.18617943241541787   0.637669698277504   0.4633804511919747   0.23037570334719007   0.34949291183722797   0.6491619401257368   0.623372682385516   0.8375011738780938   0.8082105342717611   0.7794486622550054   0.9594931206246914   0.8383063576221754   0.9467782196370653   0.6501958509685394   0.46822156955450095   0.7375783719500888   0.3970825712219472
0.7800309932874746   0.11432267922000196   0.00403520950687079   0.7451647350909066   0.6523895874550943   0.283133047582441   0.5483931405264618   0.5589853026754887   0.014719889177590359   0.8197525963904664   0.3180174371792717   0.20949239083826085   0.36555794905185357   0.19637991400495036   0.48051626330117797   0.40128185656649973   0.5861092867968482   0.23688679338025892   0.6422099056790026   0.45450363692943446   0.9359134358283088   0.768665223825758   0.9046315337289138   0.05742106570748726   0.15588244254083414   0.654342544605756   0.9005963242220429   0.3122563306165806   0.5034928550857397   0.371209497023315   0.35220318369558123   0.7532710279410918   0.4887729659081494   0.5514569006328487   0.03418574651630951   0.5437786371028309   0.12321501685629585   0.3550769866278983   0.5536694832151315   0.14249678053633127   0.5371057300594477   0.11819019324763937   0.9114595775361289   0.6879931436068968   0.601192294231139   0.3495249694218814   0.006828043807215163   0.6305720778994096   0.44530985169030485   0.6951824248161254   0.10623171958517218   0.31831574728282896   0.9418169966045651   0.32397292779281034   0.754028535889591   0.5650447193417372   0.4530440306964157   0.7725160271599617   0.7198427893732815   0.021266082238906168   0.32982901384011987   0.4174390405320634   0.16617330615814993   0.878769301702575
0.7927232837806721   0.299248847284424   0.254713728622021   0.19077615809567808   0.19153098954953315   0.9497238778625426   0.24788568481480583   0.5602040801962686   0.7462211378592284   0.25454145304641734   0.14165396522963367   0.24188833291343956   0.8044041412546633   0.930568525253607   0.3876254293400427   0.6768436135717024   0.35136011055824756   0.15805249809364533   0.6677826399667612   0.6555775313327963   0.021531096718127727   0.7406134575615819   0.5016093338086113   0.7768082296302213   0.2288078129374556   0.44136461027715795   0.24689560518659032   0.5860320715345433   0.03727682338792244   0.4916407324146153   0.9990099203717845   0.025827991338274747   0.2910556855286941   0.23709927936819797   0.8573559551421508   0.7839396584248352   0.48665154427403085   0.30653075411459096   0.4697305258021081   0.10709604485313277   0.13529143371578325   0.14847825602094564   0.8019478858353469   0.4515185135203365   0.11376033699765555   0.4078647984593637   0.3003385520267356   0.6747102838901152   0.8849525240602   0.9665001881822057   0.05344294684014529   0.08867821235557193   0.8476757006722775   0.4748594557675905   0.05443302646836081   0.06285022101729719   0.5566200151435834   0.23776017639939248   0.19707707132621   0.278910562592462   0.06996847086955256   0.9312294222848015   0.7273465455241018   0.1718145177393292
0.9346770371537693   0.7827511662638559   0.9253986596887549   0.7202960042189926   0.8209167001561137   0.3748863678044922   0.6250601076620194   0.045585720328877484   0.9359641760959139   0.4083861796222864   0.5716171608218741   0.9569075079733056   0.08828847542363633   0.9335267238546959   0.5171841343535133   0.8940572869560084   0.5316684602800529   0.6957665474553034   0.32010706302730324   0.6151467243635463   0.4616999894105004   0.764537125170502   0.5927605175032015   0.4433322066242172   0.5270229522567311   0.9817859589066461   0.6673618578144465   0.7230362024052245   0.7061062521006173   0.6068995911021539   0.04230175015242712   0.6774504820763471   0.7701420760047035   0.19851341147986745   0.47068458933055307   0.7205429741030415   0.6818536005810671   0.2649866876251715   0.9535004549770398   0.8264856871470331   0.15018514030101426   0.569220140169868   0.6333933919497365   0.21133896278348668   0.6884851508905139   0.8046830149993661   0.040632874446535135   0.7680067561592695   0.1614621986337828   0.82289705609272   0.37327101663208867   0.044970553754045024   0.4553559465331655   0.2159974649905661   0.3309692664796616   0.367520071677698   0.6852138705284619   0.017484053510698646   0.8602846771491085   0.6469770975746566   0.0033602699473948084   0.7524973658855272   0.9067842221720687   0.8204914104276235
0.8531751296463805   0.18327722571565913   0.2733908302223321   0.6091524476441368   0.16468997875586666   0.37859421071629307   0.232757955775797   0.8411456914848673   0.0032277801220838374   0.555697154623573   0.8594869391437083   0.7961751377308223   0.5478718335889183   0.33969968963300695   0.5285176726640468   0.42865506605312426   0.8626579630604564   0.3222156361223083   0.6682329955149383   0.7816779684784677   0.8592976931130616   0.5697182702367811   0.7614487733428695   0.9611865580508442   0.006122563466680992   0.386441044521122   0.48805794312053746   0.35203411040670735   0.8414325847108144   0.00784683380482897   0.25529998734474046   0.5108884189218401   0.8382048045887305   0.4521496791812559   0.39581304820103214   0.7147132811910178   0.29033297099981215   0.11244998954824899   0.8672953755369853   0.2860582151378936   0.4276750079393558   0.7902343534259407   0.19906238002204707   0.5043802466594259   0.5683773148262943   0.22051608318915955   0.4376136066791775   0.5431936886085817   0.5622547513596132   0.8340750386680376   0.9495556635586401   0.1911595782018744   0.720822166648799   0.8262282048632086   0.6942556762138996   0.6802711592800343   0.8826173620600685   0.37407852568195266   0.2984426280128675   0.9655578780890165   0.5922843910602563   0.2616285361337037   0.4311472524758821   0.6794996629511229
0.16460938312090048   0.47139418270776295   0.23208487245383505   0.17511941629169697   0.5962320682946062   0.2508780995186034   0.7944712657746575   0.6319257276831152   0.03397731693499293   0.41680306085056584   0.8449156022160176   0.4407661494812408   0.313155150286194   0.5905748559873573   0.15065992600211797   0.7604949902012065   0.43053778822612554   0.21649633030540463   0.8522172979892505   0.79493711211219   0.8382533971658692   0.954867794171701   0.4210700455133684   0.1154374491610671   0.6736440140449688   0.483473611463938   0.18898517305953333   0.9403180328693701   0.07741194575036259   0.23259551194533462   0.3945139072848758   0.30839230518625493   0.04343462881536965   0.8157924510947687   0.5495983050688582   0.8676261557050141   0.7302794785291756   0.2252175951074115   0.39893837906674023   0.1071311655038076   0.2997416903030501   0.008721264802006854   0.5467210810774897   0.3121940533916176   0.4614882931371808   0.05385347063030589   0.12565103556412133   0.19675660423055047   0.787844279092212   0.5703798591663679   0.9366658625045879   0.25643857136118037   0.7104323333418494   0.3377843472210333   0.5421519552197122   0.9480462661749254   0.6669977045264798   0.5219918961262645   0.992553650150854   0.08042011046991134   0.9367182259973041   0.29677430101885305   0.5936152710841138   0.9732889449661037
0.636976535694254   0.2880530362168462   0.046894190006624065   0.6610948915744862   0.17548824255707324   0.2341995655865403   0.9212431544425027   0.4643382873439357   0.3876439634648612   0.6638197064201724   0.9845772919379148   0.20789971598275536   0.6772116301230118   0.3260353591991391   0.44242533671820256   0.25985344980782993   0.010213925596531911   0.8040434630728747   0.44987168656734855   0.17943333933791858   0.07349569959922775   0.5072691620540216   0.8562564154832348   0.20614439437181484   0.4365191639049737   0.21921612583717542   0.8093622254766107   0.5450495027973287   0.26103092134790046   0.9850165602506351   0.888119071034108   0.08071121545339298   0.8733869578830393   0.32119685383046276   0.9035417790961932   0.8728114994706376   0.19617532776002755   0.9951614946313236   0.46111644237799065   0.6129580496628076   0.18596140216349563   0.19111803155844898   0.011244755810642066   0.4335247103248891   0.1124657025642679   0.6838488695044274   0.15498834032740727   0.22738031595307429   0.6759465386592942   0.46463274366725194   0.34562611485079653   0.6823308131557456   0.41491561731139376   0.4796161834166168   0.45750704381668855   0.6016195977023526   0.5415286594283545   0.1584193295861541   0.5539652647204953   0.728808098231715   0.34535333166832693   0.16325783495483048   0.09284882234250473   0.11585004856890731
0.15939192950483128   0.9721398033963815   0.08160406653186267   0.6823253382440182   0.046926226940563386   0.28829093389195415   0.9266157262044554   0.4549450222909439   0.3709796882812692   0.8236581902247022   0.5809896113536589   0.7726142091351983   0.9560640709698754   0.34404200680808533   0.12348256753697028   0.1709946114328457   0.41453541154152096   0.18562267722193126   0.569517302816475   0.44218651320113067   0.06918207987319407   0.02236484226710078   0.4766684804739702   0.3263364646322234   0.9097901503683627   0.05022503887071926   0.3950644139421075   0.6440111263882051   0.8628639234277994   0.7619341049787651   0.46844868773765214   0.18906610409726124   0.49188423514653024   0.9382759147540629   0.8874590763839932   0.4164518949620629   0.5358201641766548   0.5942339079459776   0.763976508847023   0.24545728352921725   0.1212847526351338   0.4086112307240463   0.1944592060305481   0.8032707703280866   0.05210267276193974   0.38624638845694553   0.7177907255565779   0.4769343056958632   0.14231252239357695   0.33602134958622626   0.3227263116144704   0.832923179307658   0.27944859896577756   0.5740872446074612   0.8542776238768183   0.6438570752103968   0.7875643638192473   0.6358113298533982   0.966818547492825   0.2274051802483339   0.25174419964259254   0.04157742190742062   0.202842038645802   0.9819478967191166
0.13045944700745873   0.6329661911833743   0.008382832615253901   0.17867712639103006   0.078356774245519   0.24671980272642877   0.290592107058676   0.7017428206951668   0.9360442518519421   0.9106984531402025   0.9678657954442056   0.8688196413875088   0.6565956528861645   0.33661120853274135   0.11358817156738736   0.224962566177112   0.8690312890669172   0.7007998786793431   0.14676962407456237   0.9975573859287781   0.6172870894243246   0.6592224567719225   0.9439275854287604   0.01560948920966146   0.4868276424168659   0.026256265588548218   0.9355447528135065   0.8369323628186314   0.40847086817134687   0.7795364628621194   0.6449526457548305   0.13518954212346454   0.47242661631940486   0.8688380097219169   0.6770868503106249   0.26636990073595573   0.8158309634332404   0.5322268011891755   0.5634986787432376   0.041407334558843746   0.9467996743663232   0.8314269225098324   0.41672905466867516   0.043849948630065645   0.32951258494199853   0.1722044657379099   0.47280146923991473   0.028240459420404183   0.8426849425251326   0.14594820014936166   0.5372567164264083   0.19130809660177278   0.43421407435378573   0.36641173728724225   0.8923040706715778   0.05611855447830825   0.9617874580343809   0.4975737275653253   0.2152172203609529   0.7897486537423525   0.14595649460114057   0.9653469263761497   0.6517185416177154   0.7483413191835088
0.19915682023481743   0.1339200038663173   0.23498948694904026   0.7044913705534431   0.8696442352928189   0.9617155381284074   0.7621880177091255   0.6762509111330389   0.026959292767686265   0.8157673379790458   0.22493130128271724   0.48494281453126614   0.5927452184139005   0.4493556006918035   0.33262723061113947   0.4288242600529579   0.6309577603795196   0.9517818731264782   0.11741001025018657   0.6390756063106053   0.48500126577837904   0.9864349467503285   0.4656914686324712   0.8907342871270966   0.28584444554356164   0.8525149428840112   0.23070198168343092   0.1862429165736535   0.4162002102507427   0.8907994047556037   0.46851396397430545   0.5099920054406145   0.38924091748305645   0.07503206677655799   0.24358266269158818   0.025049190909348405   0.796495699069156   0.6256764660847545   0.9109554320804487   0.5962249308563905   0.16553793868963634   0.6738945929582763   0.7935454218302621   0.9571493245457852   0.6805366729112573   0.6874596462079477   0.327853953197791   0.06641503741868851   0.39469222736769566   0.8349447033239366   0.09715197151436003   0.880172120845035   0.9784920171169529   0.9441452985683328   0.6286380075400546   0.3701801154044205   0.5892510996338964   0.8691132317917748   0.38505534484846643   0.34513092449507204   0.7927554005647405   0.24343676570702036   0.4740999127680177   0.7489059936386815
0.6272174618751042   0.5695421727487441   0.6805544909377556   0.7917566690928964   0.9466807889638469   0.8820825265407963   0.3527005377399646   0.725341631674208   0.5519885615961513   0.04713782321685974   0.25554856622560457   0.8451695108291729   0.5734965444791983   0.1029925246485269   0.62691055868555   0.47498939542475244   0.9842454448453019   0.23387929285675205   0.24185521383708358   0.1298584709296804   0.1914900442805613   0.9904425271497317   0.7677553010690659   0.38095247729099885   0.5642725824054571   0.4209003544009876   0.0872008101313103   0.5891958081981025   0.6175917934416102   0.5388178278601913   0.7345002723913457   0.8638541765238945   0.06560323184545898   0.4916800046433315   0.4789517061657411   0.01868466569472162   0.4921066873662607   0.38868747999480463   0.8520411474801911   0.5436952702699692   0.5078612425209589   0.15480818713805256   0.6101859336431075   0.4138367993402888   0.31637119824039756   0.16436565998832087   0.8424306325740416   0.032884322049289906   0.7520986158349404   0.7434653055873333   0.7552298224427313   0.44368851385118746   0.13450682239333026   0.204647477727142   0.02072955005138566   0.579834337327293   0.06890359054787128   0.7129674730838105   0.5417778438856445   0.5611496716325713   0.5767969031816106   0.32427999308900585   0.6897366964054534   0.017454401362602154
0.06893566066065171   0.1694718059509533   0.07955076276234593   0.6036176020223134   0.7525644624202541   0.005106145962632426   0.23712013018830427   0.5707332799730235   0.0004658465853136643   0.26164084037529917   0.48189030774557295   0.12704476612183602   0.8659590241919835   0.05699336264815715   0.4611607576941873   0.5472104287945431   0.7970554336441121   0.34402588956434665   0.9193829138085428   0.9860607571619717   0.22025853046250157   0.01974589647534081   0.22964621740308927   0.9686063557993696   0.15132286980184986   0.8502740905243875   0.15009545464074334   0.3649887537770562   0.39875840738159574   0.8451679445617551   0.912975324452439   0.7942554738040327   0.39829256079628206   0.5835271041864559   0.4310850167068661   0.6672107076821967   0.5323335366042986   0.5265337415382988   0.9699242590126789   0.12000027888765365   0.7352781029601865   0.1825078519739521   0.05054134520413611   0.1339395217256819   0.5150195724976849   0.1627619554986113   0.8208951278010469   0.1653331659263123   0.3636967026958351   0.31248786497422376   0.6707996731603035   0.8003444121492561   0.9649382953142394   0.46731992041246867   0.7578243487078645   0.006088938345223391   0.5666457345179573   0.8837928162260128   0.32673933200099836   0.3388782306630267   0.03431219791365866   0.35725907468771395   0.35681507298831955   0.21887795177537303
0.29903409495347216   0.17475122271376187   0.30627372778418344   0.08493843004969111   0.7840145224557872   0.01198926721515055   0.4853785999831366   0.9196052641233788   0.4203178197599521   0.6995014022409267   0.8145789268228331   0.11926085197412267   0.4553795244457127   0.23218148182845808   0.05675457811496858   0.11317191362889928   0.8887337899277554   0.3483886656024453   0.7300152461139702   0.7742936829658726   0.8544215920140967   0.9911295909147313   0.3732001731256507   0.5554157311904996   0.5553874970606246   0.8163783682009695   0.06692644534146726   0.4704773011408085   0.7713729746048374   0.804389100985819   0.5815478453583307   0.5508720370174297   0.3510551548448853   0.10488769874489218   0.7669689185354976   0.43161118504330703   0.8956756303991725   0.8727062169164341   0.710214340420529   0.31843927141440775   0.006941840471417149   0.5243175513139888   0.9801990943065588   0.5441455884485351   0.15252024845732037   0.5331879603992574   0.6069989211809081   0.9887298572580355   0.5971327513966957   0.716809592198288   0.5400724758394408   0.5182525561172271   0.8257597767918583   0.912420491212469   0.9585246304811101   0.9673805190997974   0.47470462194697305   0.8075327924675768   0.19155571194561255   0.5357693340564904   0.5790289915478005   0.9348265755511427   0.4813413715250835   0.21733006264208263
0.5720871510763833   0.4105090242371539   0.5011422772185247   0.6731844741935475   0.41956690261906293   0.8773210638378964   0.8941433560376165   0.6844546169355119   0.8224341512223672   0.16051147163960855   0.3540708801981756   0.16620206081828487   0.9966743744305088   0.24809098042713953   0.3955462497170654   0.1988215417184875   0.5219697524835357   0.4405581879595627   0.20399053777145287   0.6630522076619971   0.9429407609357353   0.50573161240842   0.7226491662463693   0.44572214501991453   0.370853609859352   0.09522258817126608   0.2215068890278447   0.772537670826367   0.9512867072402891   0.2179015243333696   0.3273635329902282   0.08808305389085508   0.12885255601792187   0.05739005269376106   0.9732926527920526   0.9218809930725702   0.13217818158741307   0.8092990722666216   0.5777464030749871   0.7230594513540827   0.6102084291038773   0.3687408843070588   0.3737558653035342   0.060007243692085564   0.667267668168142   0.8630092718986387   0.6511066990571649   0.6142850986721711   0.29641405830879003   0.7677866837273727   0.42959981002932013   0.841747427845804   0.34512735106850095   0.5498851593940032   0.10223627703909195   0.7536643739549489   0.2162747950505791   0.49249510670024205   0.1289436242470394   0.8317833808823787   0.08409661346316602   0.6831960344336205   0.5511972211720523   0.10872392952829603
0.4738881843592887   0.3144551501265617   0.17744135586851809   0.04871668583621047   0.8066205161911467   0.4514458782279229   0.5263346568113533   0.4344315871640394   0.5102064578823567   0.6836591945005502   0.09673484678203309   0.5926841593182354   0.16507910681385576   0.13377403510654712   0.9944985697429412   0.8390197853632865   0.9488043117632767   0.6412789284063051   0.8655549454959017   0.007236404480907732   0.8647076983001106   0.9580828939726845   0.31435772432384945   0.8985124749526117   0.3908195139408219   0.6436277438461228   0.13691636845533137   0.8497957891164012   0.5841989977496752   0.1921818656181998   0.6105817116439781   0.4153642019523618   0.07399253986731848   0.5085226711176496   0.513846864861945   0.8226800426341264   0.9089134330534627   0.3747486360111025   0.5193482951190039   0.9836602572708399   0.960109121290186   0.7334697076047975   0.6537933496231022   0.9764238527899322   0.09540142299007533   0.7753868136321129   0.3394356252992527   0.0779113778373205   0.7045819090492533   0.13175906978599017   0.20251925684392136   0.22811558872091928   0.12038291129957816   0.9395772041677903   0.5919375451999432   0.8127513867685575   0.04639037143225968   0.43105453305014074   0.07809068033799821   0.9900713441344311   0.137476938378797   0.056305897039038294   0.5587423852189943   0.006411086863591136
0.17736781708861096   0.32283618943424086   0.9049490355958921   0.029987234073658938   0.08196639409853564   0.5474493758021279   0.5655134102966395   0.9520758562363384   0.3773844850492823   0.41569030601613777   0.36299415345271807   0.7239602675154192   0.2570015737497041   0.47611310184834743   0.7710566082527749   0.9112088807468617   0.21061120231744443   0.04505856879820666   0.6929659279147766   0.9211375366124306   0.07313426393864744   0.9887526717591684   0.1342235426957823   0.9147264497488395   0.8957664468500365   0.6659164823249275   0.22927450709989014   0.8847392156751805   0.8138000527515008   0.11846710652279956   0.6637610968032507   0.9326633594388422   0.43641556770221857   0.7027768005066618   0.3007669433505326   0.20870309192342296   0.17941399395251448   0.22666369865831434   0.5297103350977578   0.2974942111765613   0.96880279163507   0.18160512986010768   0.8367444071829812   0.37635667456413063   0.8956685276964226   0.19285245810093932   0.7025208644871989   0.46163022481529115   0.9999020808463861   0.5269359757760118   0.4732463573873087   0.5768910091401106   0.1861020280948853   0.4084688692532123   0.809485260584058   0.6442276497012684   0.7496864603926667   0.7056920687465505   0.5087183172335255   0.4355245577778455   0.5702724664401523   0.4790283700882362   0.9790079821357677   0.13803034660128424
0.6014696748050822   0.2974232402281285   0.14226357495278652   0.7616736720371536   0.7058011471086596   0.10457078212718915   0.4397427104655877   0.3000434472218625   0.7058990662622735   0.5776348063511774   0.966496353078279   0.7231524380817519   0.5197970381673882   0.16916593709796504   0.157011092494221   0.07892478838048347   0.7701105777747215   0.4634738683514145   0.6482927752606955   0.643400230602638   0.19983811133456922   0.9844454982631784   0.669284793124928   0.5053698840013537   0.598368436529487   0.6870222580350499   0.5270212181721413   0.7436962119642001   0.8925672894208274   0.5824514759078607   0.08727850770655365   0.4436527647423376   0.18666822315855391   0.004816669556683438   0.12078215462827466   0.7205003266605857   0.6668711849911657   0.8356507324587183   0.9637710621340537   0.6415755382801023   0.8967606072164442   0.3721768641073039   0.3154782868733581   0.9981753076774643   0.696922495881875   0.3877313658441255   0.6461934937484303   0.4928054236761105   0.098554059352388   0.7007091078090756   0.11917227557628887   0.7491092117119104   0.2059867699315606   0.11825763190121484   0.03189376786973521   0.3054564469695728   0.019318546773006654   0.1134409623445314   0.9111116132414605   0.584956120308987   0.35244736178184094   0.277790229885813   0.9473405511074069   0.9433805820288849
0.4556867545653967   0.9056133657785091   0.6318622642340488   0.9452052743514205   0.7587642586835217   0.5178819999343837   0.9856687704856185   0.45239985067531   0.6602101993311337   0.8171728921253081   0.8664964949093297   0.7032906389633996   0.45422342939957305   0.6989152602240932   0.8346027270395945   0.39783419199382686   0.4349048826265664   0.5854742978795618   0.9234911137981339   0.8128780716848397   0.0824575208447255   0.3076840679937488   0.976150562690727   0.869497489655955   0.6267707662793288   0.40207070221523966   0.3442882984566783   0.9242922153045343   0.8680065075958072   0.884188702280856   0.3586195279710598   0.47189236462922435   0.20779630826467352   0.06701581015554799   0.4921230330617301   0.7686017256658247   0.7535728788651004   0.3681005499314548   0.6575203060221357   0.37076753367199783   0.318667996238534   0.782626252051893   0.7340291922240018   0.557889461987158   0.23621047539380852   0.47494218405814415   0.7578786295332748   0.6883919723312031   0.6094397091144796   0.07287148184290447   0.4135903310765965   0.7640997570266688   0.7414332015186725   0.18868277956204843   0.05497080310553673   0.2922073923974444   0.533636893253999   0.12166696940650044   0.5628477700438066   0.5236056667316198   0.7800640143888986   0.7535664194750457   0.905327464021671   0.1528381330596219
0.4613960181503646   0.9709401674231527   0.1712982717976691   0.5949486710724639   0.22518554275655608   0.49599798336500855   0.4134196422643943   0.9065566987412607   0.6157458336420764   0.42312650152210407   0.9998293111877978   0.14245694171459194   0.8743126321234039   0.23444372196005564   0.9448585080822611   0.8502495493171475   0.3406757388694049   0.1127767525535552   0.3820107380384545   0.3266438825855278   0.5606117244805063   0.3592103330785095   0.47668327401678356   0.17380574952590588   0.0992157063301417   0.3882701656553568   0.30538500221911447   0.578857078453442   0.8740301635735857   0.8922721822903483   0.8919653599547201   0.6723003797121814   0.25828432993150924   0.4691456807682442   0.8921360487669223   0.5298434379975894   0.38397169780810536   0.23470195880818856   0.9472775406846612   0.6795938886804419   0.04329595893870048   0.12192520625463335   0.5652668026462068   0.3529500060949141   0.4826842344581942   0.7627148731761239   0.08858352862942316   0.17914425656900826   0.3834685281280525   0.374444707520767   0.7831985264103087   0.6002871781155662   0.5094383645544669   0.4821725252304187   0.8912331664555886   0.9279867984033848   0.2511540346229576   0.013026844462174513   0.9990971176886663   0.39814336040579545   0.8671823368148522   0.7783248856539859   0.051819577004005045   0.7185494717253536
0.8238863778761518   0.6563996793993526   0.4865527743577983   0.3655994656304395   0.34120214341795757   0.8936848062232288   0.39796924572837516   0.18645520906143123   0.9577336152899051   0.5192400987024618   0.6147707193180665   0.586168030945865   0.44829525073543824   0.037067573472043105   0.7235375528624779   0.6581812325424802   0.19714121611248067   0.02404072900986859   0.7244404351738116   0.26003787213668467   0.3299588792976284   0.24571584335588262   0.6726208581698065   0.5414884004113311   0.5060725014214766   0.58931616395653   0.18606808381200826   0.17588893478089163   0.16487035800351904   0.6956313577333012   0.7880988380836331   0.9894337257194604   0.20713674271361393   0.1763912590308394   0.17332811876556667   0.40326569477359536   0.7588414919781756   0.1393236855587963   0.4497905659030888   0.7450844622311152   0.561700275865695   0.1152829565489277   0.7253501307292771   0.4850465900944306   0.23174139656806658   0.869567113193045   0.05272927255947059   0.9435581896830995   0.7256688951465899   0.28025094923651506   0.8666611887474623   0.7676692549022078   0.5607985371430709   0.5846195915032139   0.07856235066382923   0.7782355291827475   0.353661794429457   0.40822833247237444   0.9052342318982626   0.3749698344091521   0.5948203024512814   0.2689046469135782   0.4554436659951738   0.6298853721780369
0.03312002658558636   0.15362169036465045   0.7300935352658966   0.1448387820836063   0.8013786300175197   0.28405457717160537   0.677364262706426   0.2012805924005068   0.07570973487092982   0.003803627935090307   0.8107030739589637   0.43361133749829894   0.5149111977278589   0.41918403643187646   0.7321407232951345   0.6553758083155514   0.1612494032984019   0.010955703959501982   0.8269064913968719   0.2804059739063994   0.5664291008471205   0.7420510570459238   0.3714628254016981   0.6505206017283626   0.5333090742615342   0.5884293666812733   0.6413692901358015   0.5056818196447562   0.7319304442440144   0.30437478950966795   0.9640050274293754   0.30440122724424945   0.6562207093730846   0.3005711615745777   0.15330195347041176   0.8707898897459505   0.14130951164522568   0.8813871251427012   0.42116123017527723   0.21541408143039903   0.9800601083468238   0.8704314211831993   0.5942547387784053   0.9350081075239997   0.4136310074997033   0.12838036413727544   0.2227919133767072   0.2844875057956371   0.8803219332381691   0.5399509974560021   0.5814226232409057   0.7788056861508809   0.14839148899415466   0.2355762079463341   0.6174175958115302   0.4744044589066314   0.4921707796210701   0.9350050463717564   0.4641156423411185   0.6036145691606809   0.35086126797584444   0.05361792122905521   0.04295441216584125   0.38820048773028193
0.3708011596290206   0.18318650004585596   0.4486996733874359   0.4531923802062823   0.9571701521293173   0.05480613590858054   0.2259077600107287   0.16870487441064516   0.0768482188911483   0.5148551384525785   0.644485136769823   0.3898991882597643   0.9284567298969937   0.27927893050624436   0.027067540958292745   0.9154947293531329   0.43628595027592354   0.34427388413448795   0.5629518986171742   0.31188016019245196   0.08542468230007912   0.2906559629054327   0.519997486451333   0.9236796724621701   0.7146235226710584   0.10746946285957677   0.07129781306389708   0.47048729225588776   0.7574533705417411   0.05266332695099622   0.8453900530531684   0.3017824178452426   0.6806051516505928   0.5378081884984177   0.2009049162833454   0.9118832295854783   0.7521484217535992   0.25852925799217336   0.17383737532505264   0.9963885002323455   0.31586247147767565   0.9142553738576854   0.6108854767078784   0.6845083400398935   0.23043778917759652   0.6235994109522527   0.09088799025654541   0.7608286675777235   0.515814266506538   0.5161299480926759   0.01959017719264832   0.2903413753218357   0.7583608959647969   0.4634666211416797   0.17420012413947994   0.9885589574765931   0.07775574431420415   0.925658432643262   0.9732952078561345   0.07667572789111472   0.325607322560605   0.6671291746510886   0.7994578325310819   0.08028722765876928
0.009744851082929367   0.7528738007934032   0.18857235582320347   0.3957788876188758   0.7793070619053328   0.12927438984115044   0.09768436556665808   0.6349502200411523   0.26349279539879483   0.6131444417484745   0.07809418837400976   0.3446088447193167   0.5051318994339978   0.14967782060679483   0.9038940642345298   0.35604988724272363   0.4273761551197937   0.22401938796353288   0.9305988563783952   0.2793741593516089   0.10176883255918871   0.5568902133124443   0.13114102384731338   0.19908693169283964   0.09202398147625934   0.8040164125190411   0.9425686680241099   0.8033080440739638   0.3127169195709265   0.6747420226778907   0.8448843024574518   0.1683578240328115   0.04922412417213169   0.06159758092941616   0.7667901140834421   0.8237489793134948   0.5440922247381338   0.9119197603226213   0.8628960498489122   0.46769909207077115   0.11671606961834012   0.6879003723590884   0.932297193470517   0.18832493271916226   0.014947237059151406   0.13101015904664415   0.8011561696232036   0.9892380010263226   0.922923255582892   0.326993746527603   0.8585875015990937   0.18592995695235878   0.6102063360119656   0.6522517238497123   0.013703199141641855   0.017572132919547297   0.5609822118398339   0.5906541429202962   0.24691308505819978   0.19382315360605248   0.01688998710170004   0.6787343825976748   0.38401703520928754   0.7261240615352813
0.90017391748336   0.9908340102385864   0.4517198417387706   0.537799128816119   0.8852266804242085   0.8598238511919423   0.650563672115567   0.5485611277897965   0.9623034248413165   0.5328301046643392   0.7919761705164733   0.3626311708374377   0.35209708882935087   0.8805783808146269   0.7782729713748315   0.34505903791789033   0.791114876989517   0.28992423789433075   0.5313598863166317   0.15123588431183788   0.774224889887817   0.6111898552966559   0.14734285110734413   0.42511182277655657   0.8740509724044571   0.6203558450580695   0.6956230093685736   0.8873126939604374   0.9888242919802486   0.7605319938661274   0.045059337253006544   0.33875156617064106   0.026520867138932105   0.2277018892017881   0.2530831667365332   0.9761203953332034   0.6744237783095812   0.3471235083871612   0.4748101953617017   0.631061357415313   0.8833089013200642   0.05719927049283045   0.94345030904507   0.4798254731034752   0.10908401143224719   0.44600941519617454   0.7961074579377259   0.054713650326918606   0.23503303902779013   0.825653570138105   0.10048444856915234   0.1674009563664811   0.24620874704754156   0.06512157627197769   0.055425111316145796   0.82864939019584   0.21968787990860947   0.8374196870701895   0.8023419445796126   0.8525289948626367   0.5452641015990283   0.4902961786830284   0.3275317492179109   0.22146763744732367
0.661955200278964   0.43309690819019797   0.38408144017284085   0.7416421643438486   0.5528711888467168   0.9870874929940234   0.587973982235115   0.6869285140169299   0.3178381498189268   0.16143392285591843   0.4874895336659626   0.5195275576504488   0.0716294027713852   0.09631234658394074   0.4320644223498168   0.6908781674546087   0.8519415228627757   0.2588926595137511   0.6297224777702042   0.838349172591972   0.3066774212637475   0.7685964808307227   0.30219072855229334   0.6168815351446484   0.6447222209847834   0.33549957264052477   0.9181092883794525   0.8752393708007998   0.09185103213806654   0.34841207964650134   0.33013530614433756   0.1883108567838699   0.7740128823191398   0.18697815679058294   0.8426457724783749   0.6687832991334212   0.7023834795477546   0.0906658102066422   0.4105813501285581   0.9779051316788124   0.8504419566849789   0.831773150692891   0.7808588723583539   0.13955595908684043   0.5437645354212314   0.06317666986216831   0.47866814380606054   0.5226744239421921   0.8990423144364479   0.7276770972216435   0.560558855426608   0.6474350531413923   0.8071912822983814   0.3792650175751422   0.23042354928227046   0.4591241963575224   0.03317839997924161   0.19228686078455923   0.3877777768038955   0.7903408972241013   0.330794920431487   0.10162105057791704   0.9771964266753373   0.8124357655452888
0.48035296374650815   0.269847899885026   0.19633755431698344   0.6728798064584484   0.9365884283252768   0.20667123002285767   0.7176694105109229   0.15020538251625626   0.03754611388882885   0.4789941328012141   0.15711055508431485   0.502770329374864   0.23035483159044745   0.09972911522607196   0.9266870058020443   0.0436461330173416   0.19717643161120585   0.9074422544415127   0.5389092289981489   0.2533052357932404   0.8663815111797188   0.8058212038635957   0.5617128023228115   0.4408694702479516   0.3860285474332107   0.5359733039785697   0.36537524800582805   0.7679896637895032   0.44944011910793386   0.32930207395571204   0.6477058374949052   0.617784281273247   0.411894005219105   0.8503079411544979   0.49059528241059036   0.11501395189838301   0.18153917362865757   0.750578825928426   0.563908276608546   0.0713678188810414   0.9843627420174518   0.8431365714869132   0.024999047610397118   0.818062583087801   0.11798123083773289   0.03731536762331756   0.4632862452875856   0.37719311283984946   0.7319526834045222   0.5013420636447479   0.09791099728175755   0.6092034490503463   0.28251256429658833   0.17203998968903578   0.4502051597868524   0.9914191677770993   0.8706185590774833   0.32173204853453785   0.959609877376262   0.8764052158787162   0.6890793854488257   0.5711532226061119   0.39570160076771604   0.8050373969976748
0.704716643431374   0.7280166511191987   0.3707025531573189   0.9869748139098738   0.5867354125936411   0.6907012834958811   0.9074163078697333   0.6097817010700244   0.8547827291891189   0.18935921985113324   0.8095053105879757   0.000578252019678101   0.5722701648925306   0.01731923016209745   0.3593001508011234   0.009159084242578835   0.7016516058150473   0.6955871816275596   0.39969027342486135   0.13275386836386258   0.012572220366221522   0.12443395902144772   0.00398867265714535   0.32771647136618776   0.3078555769348475   0.3964173079022491   0.6332861194998265   0.3407416574563139   0.7211201643412064   0.705716024406368   0.7258698116300931   0.7309599563862896   0.8663374351520875   0.5163568045552348   0.9163645010421174   0.7303817043666114   0.29406727025955687   0.49903757439313734   0.557064350240994   0.7212226201240326   0.5924156644445097   0.8034503927655777   0.15737407681613264   0.5884687517601701   0.5798434440782881   0.67901643374413   0.1533854041589873   0.26075228039398235   0.2719878671434406   0.2825991258418809   0.5200992846591609   0.9200106229376684   0.5508677028022342   0.5768831014355129   0.7942294730290677   0.18905066655137884   0.6845302676501468   0.060526296880278115   0.8778649719869503   0.4586689621847673   0.39046299739058987   0.5614887224871408   0.32080062174595625   0.7374463420607347
0.7980473329460803   0.758038329721563   0.16342654492982364   0.14897759030056462   0.21820388886779218   0.07902189597743303   0.010041140770836336   0.8882253099065823   0.9462160217243516   0.7964227701355521   0.48994185611167546   0.9682146869689139   0.39534831892211736   0.21953966870003921   0.6957123830826077   0.7791640204175351   0.7108180512719706   0.1590133718197611   0.8178474110956575   0.3204950582327677   0.32035505388138075   0.5975246493326203   0.4970467893497012   0.583048716172033   0.5223077209353004   0.8394863196110572   0.3336202444198776   0.4340711258714684   0.30410383206750824   0.7604644236336242   0.32357910364904124   0.5458458159648861   0.3578878103431567   0.9640416534980721   0.8336372475373658   0.5776311289959722   0.9625394914210393   0.7445019847980329   0.137924864454758   0.7984671085784372   0.2517214401490687   0.5854886129782718   0.3200774533591005   0.4779720503456695   0.931366386267688   0.9879639636456515   0.8230306640093993   0.8949233341736365   0.40905866533238755   0.1484776440345942   0.4894104195895217   0.46085220830216805   0.10495483326487927   0.38801322040096997   0.16583131594048048   0.915006392337282   0.7470670229217226   0.42397156690289783   0.3321940684031147   0.3373752633413098   0.7845275315006833   0.679469582104865   0.19426920394835673   0.5389081547628727
0.5328060913516146   0.09398096912659315   0.8741917505892562   0.06093610441720317   0.6014397050839266   0.10601700548094166   0.051161086579856956   0.16601277024356673   0.19238103975153908   0.9575393614463474   0.5617506669903353   0.7051605619413986   0.08742620648665983   0.5695261410453775   0.39591935104985476   0.7901541696041167   0.3403591835649372   0.1455545741424796   0.06372528264674004   0.45277890626280687   0.555831652064254   0.46608499203761466   0.8694560786983833   0.9138707514999342   0.023025560712639358   0.3721040229110215   0.995264328109127   0.852934647082731   0.42158585562871276   0.26608701743007984   0.94410324152927   0.6869218768391644   0.22920481587717365   0.3085476559837324   0.38235257453893484   0.9817613148977657   0.14177860939051382   0.739021514938355   0.9864332234890801   0.19160714529364903   0.8014194258255766   0.5934669407958754   0.9227079408423401   0.7388282390308422   0.24558777376132265   0.1273819487582607   0.05325186214395673   0.8249574875309079   0.2225622130486833   0.7552779258472392   0.057987534034829674   0.9720228404481769   0.8009763574199705   0.48919090841715934   0.11388429250555956   0.28510096360901255   0.5717715415427969   0.18064325243342694   0.7315317179666248   0.30333964871124686   0.42999293215228307   0.441621737495072   0.7450984944775446   0.1117325034175978
0.6285735063267065   0.8481547966991966   0.8223905536352045   0.3729042643867556   0.3829857325653838   0.7207728479409359   0.7691386914912478   0.5479467768558477   0.16042351951670056   0.9654949220936967   0.7111511574564181   0.5759239364076708   0.35944716209673   0.4763040136765374   0.5972668649508586   0.2908229727986583   0.7876756205539331   0.29566076124311047   0.8657351469842339   0.9874833240874115   0.35768268840165   0.8540390237480385   0.12063665250668928   0.8757508206698137   0.7291091820749436   0.005884227048841856   0.29824609887148473   0.5028465562830581   0.34612344950955976   0.28511137910790596   0.5291074073802369   0.9548997794272103   0.18569992999285917   0.3196164570142092   0.8179562499238188   0.3789758430195395   0.8262527678961292   0.8433124433376719   0.22068938497296012   0.0881528702208812   0.038577147342196076   0.5476516820945614   0.3549542379887262   0.10066954613346973   0.680894458940546   0.6936126583465229   0.23431758548203696   0.22491872546365607   0.9517852768656024   0.687728431297681   0.9360714866105523   0.722072169180598   0.6056618273560428   0.4026170521897751   0.40696407923031536   0.7671723897533878   0.41996189736318357   0.08300059517556589   0.5890078293064966   0.38819654673384824   0.5937091294670543   0.23968815183789408   0.3683184443335365   0.30004367651296704
0.5551319821248583   0.6920364697433327   0.013364206344810267   0.1993741303794973   0.8742375231843122   0.9984238113968098   0.7790466208627733   0.9744554049158413   0.9224522463187098   0.3106953800991288   0.842975134252221   0.2523832357352432   0.3167904189626671   0.9080783279093537   0.4360110550219057   0.4852108459818555   0.8968285215994835   0.8250777327337878   0.8470032257154091   0.09701429924800722   0.3031193921324291   0.5853895808958938   0.47868478138187254   0.7969706227350402   0.7479874100075709   0.893353111152561   0.46532057503706226   0.5975964923555429   0.8737498868232585   0.8949292997557512   0.6862739541742889   0.6231410874397016   0.9512976405045488   0.5842339196566224   0.8432988199220679   0.37075785170445846   0.6345072215418817   0.6761555917472688   0.4072877649001622   0.8855470057226029   0.7376786999423982   0.851077859013481   0.5602845391847532   0.7885327064745957   0.4345593078099691   0.2656882781175873   0.08159975780288062   0.9915620837395556   0.6865718978023982   0.3723351669650262   0.6162791827658184   0.3939655913840127   0.8128220109791398   0.477405867209275   0.9300052285915293   0.770824503944311   0.861524370474591   0.8931719475526526   0.08670640866946146   0.4000666522398526   0.22701714893270927   0.21701635580538384   0.6794186437692993   0.5145196465172497
0.4893384489903111   0.3659384967919029   0.11913410458454607   0.7259869400426538   0.054779141180341974   0.10025021867431562   0.03753434678166545   0.7344248563030983   0.3682072433779437   0.7279150517092894   0.4212551640158471   0.3404592649190856   0.555385232398804   0.25050918450001436   0.4912499354243177   0.5696347609747746   0.693860861924213   0.35733723694736175   0.4045435267548563   0.16956810873492198   0.46684371299150373   0.1403208811419779   0.7251248829855571   0.6550484622176723   0.9775052640011926   0.774382384350075   0.605990778401011   0.9290615221750185   0.9227261228208506   0.6741321656757594   0.5684564316193456   0.1946366658719201   0.554518879442907   0.94621711396647   0.14720126760349841   0.8541774009528345   0.999133647044103   0.6957079294664557   0.6559513321791807   0.28454263997805984   0.30527278511989003   0.33837069251909396   0.2514078054243244   0.11497453124313789   0.8384290721283864   0.19804981137711605   0.5262829224387674   0.45992606902546557   0.8609238081271936   0.423667427027041   0.9202921440377564   0.5308645468504471   0.938197685306343   0.7495352613512816   0.35183571241841083   0.336227880978527   0.383678805863436   0.8033181473848116   0.20463444481491241   0.48205048002569256   0.384545158819333   0.10761021791835579   0.5486831126357317   0.19750784004763267
0.07927237369944296   0.7692395253992619   0.2972753072114073   0.08253330880449479   0.24084330157105666   0.5711897140221458   0.77099238477264   0.6226072397790292   0.379919493443863   0.1475222869951048   0.8507002407348836   0.09174269292858214   0.44172180813752   0.39798702564382327   0.49886452831647277   0.7555148119500551   0.05804300227408402   0.5946688782590117   0.2942300835015604   0.2734643319243626   0.673497843454751   0.4870586603406559   0.7455469708658287   0.07595649187672991   0.5942254697553081   0.7178191349413942   0.44827166365442134   0.9934231830722351   0.35338216818425144   0.1466294209192483   0.6772792788817814   0.3708159432932059   0.9734626747403885   0.9991071339241435   0.8265790381468978   0.2790732503646237   0.5317408666028685   0.6011201082803203   0.327714509830425   0.5235584384145686   0.4736978643287844   0.006451230021308526   0.03348442632886463   0.250094106490206   0.8002000208740334   0.5193925696806526   0.28793745546303595   0.1741376146134761   0.20597455111872529   0.8015734347392585   0.8396657918086147   0.18071443154124098   0.8525923829344738   0.6549440138200102   0.16238651292683326   0.8098984882480351   0.8791297081940853   0.6558368798958667   0.3358074747799355   0.5308252378834114   0.3473888415912169   0.0547167716155464   0.008092964949510482   0.007266799468842762
0.8736909772624325   0.048265541594237876   0.9746085386206459   0.7571726929786368   0.07349095638839911   0.5288729719135853   0.6866710831576099   0.5830350783651607   0.8675164052696739   0.7272995371743268   0.8470052913489953   0.40232064682391966   0.014924022335200007   0.07235552335431665   0.684618778422162   0.5924221585758845   0.13579431414111465   0.41651864345844997   0.3488113036422265   0.06159692069247321   0.7884054725498977   0.3618018718429036   0.34071833869271606   0.05433012122363044   0.9147144952874653   0.31353633024866573   0.3661098000720702   0.2971574282449937   0.8412235388990661   0.7846633583350804   0.6794387169144603   0.714122349879833   0.9737071336293923   0.0573638211607536   0.8324334255654651   0.31180170305591337   0.9587831112941922   0.985008297806437   0.14781464714330303   0.7193795444800288   0.8229887971530776   0.5684896543479869   0.7990033435010765   0.6577826237875556   0.03458332460317992   0.2066877825050834   0.45828500480836043   0.6034525025639251   0.11986882931571467   0.8931514522564177   0.09217520473629025   0.30629507431893144   0.27864529041664854   0.10848809392133728   0.4127364878218299   0.5921727244390984   0.3049381567872562   0.05112427276058368   0.5803030622563649   0.28037102138318504   0.3461550454930639   0.06611597495414671   0.43248841511306185   0.5609914769031562
0.5231662483399863   0.49762632060615974   0.6334850716119854   0.9032088531156007   0.48858292373680634   0.29093853810107634   0.17520006680362493   0.29975635055167554   0.3687140944210917   0.39778708584465866   0.08302486206733467   0.993461276232744   0.09006880400444316   0.28929899192332137   0.6702883742455047   0.4012885517936457   0.785130647217187   0.2381747191627377   0.08998531198913984   0.12091753041046065   0.438975601724123   0.172058744208591   0.6574968968760779   0.5599260535073044   0.9158093533841367   0.6744324236024313   0.024011825264092613   0.6567172003917037   0.4272264296473303   0.3834938855013549   0.8488117584604677   0.3569608498400282   0.05851233522623865   0.9857067996566963   0.765786896393133   0.3634995736072841   0.9684435312217955   0.6964078077333749   0.09549852214762829   0.9622110218136384   0.18331288400460857   0.45823308857063716   0.0055132101584884526   0.8412934914031778   0.7443372822804856   0.2861743443620462   0.34801631328241045   0.2813674378958733   0.8285279288963489   0.611741920759615   0.3240044880183179   0.6246502375041696   0.40130149924901853   0.22824803525826004   0.4751927295578502   0.26768938766414146   0.34278916402277987   0.2425412356015638   0.7094058331647172   0.9041898140568574   0.3743456328009844   0.546133427868189   0.6139073110170888   0.941978792243219
0.1910327487963758   0.0879003392975518   0.6083941008586004   0.10068530084004124   0.4466954665158902   0.8017259949355057   0.2603777875761899   0.8193178629441679   0.6181675376195414   0.1899840741758907   0.9363732995578721   0.19466762543999827   0.21686603837052282   0.9617360389176307   0.4611805700000219   0.9269782377758569   0.874076874347743   0.7191948033160669   0.7517747368353047   0.022788423718999466   0.4997312415467585   0.17306137544787792   0.1378674258182159   0.08080963147578049   0.30869849275038275   0.08516103615032611   0.5294733249596155   0.9801243306357392   0.8620030262344925   0.2834350412148205   0.26909553738342556   0.16080646769157136   0.24383548861495113   0.09345096703892979   0.33272223782555355   0.9661388422515731   0.02696945024442833   0.13171492812129912   0.8715416678255317   0.03916060447571629   0.1528925758966854   0.41252012480523226   0.11976693099022687   0.016372180756716818   0.6531613343499268   0.23945874935735437   0.981899505172011   0.9355625492809363   0.34446284159954416   0.15429771320702826   0.45242618021239545   0.9554382186451971   0.4824598153650516   0.8708626719922078   0.18333064282896988   0.7946317509536257   0.23862432675010048   0.7774117049532779   0.8506084050034164   0.8284929087020526   0.21165487650567216   0.6456967768319789   0.9790667371778847   0.7893323042263363
0.05876230060898675   0.2331766520267466   0.8592998061876579   0.7729601234696195   0.4056009662590599   0.9937179026693922   0.8774003010156469   0.8373975741886831   0.061138124659515763   0.839420189462364   0.4249741208032514   0.881959355543486   0.5786783092944642   0.9685575174701562   0.24164347797428154   0.0873276045898604   0.34005398254436364   0.19114581251687823   0.3910350729708652   0.25883469588780783   0.1283991060386915   0.5454490356848993   0.4119683357929805   0.46950239166147156   0.06963680542970474   0.3122723836581528   0.5526685296053226   0.696542268191852   0.6640358391706449   0.31855448098876055   0.6752682285896757   0.859144694003169   0.6028977145111291   0.4791342915263965   0.2502941077864243   0.9771853384596828   0.02421940521666495   0.5105767740562404   0.008650629812142728   0.8898577338698225   0.6841654226723013   0.3194309615393621   0.6176155568412776   0.6310230379820146   0.5557663166336098   0.7739819258544628   0.20564722104829708   0.16152064632054305   0.4861295112039051   0.46170954219631   0.6529786914429745   0.464978378128691   0.8220936720332602   0.14315506120754942   0.9777104628532988   0.6058336841255221   0.2191959575221311   0.6640207696811529   0.7274163550668745   0.6286483456658392   0.19497655230546618   0.15344399562491254   0.7187657252547318   0.7387906117960167
0.5108111296331649   0.8340130340855504   0.10115016841345423   0.10776757381400211   0.9550448129995551   0.06003110823108768   0.8955029473651571   0.9462469274934591   0.46891530179565   0.5983215660347777   0.24252425592218269   0.4812685493647681   0.6468216297623898   0.45516650482722826   0.2648137930688839   0.8754348652392461   0.42762567224025866   0.7911457351460754   0.5373974380020095   0.24678651957340686   0.2326491199347925   0.6377017395211628   0.8186317127472776   0.5079959077773901   0.7218379903016277   0.8036887054356124   0.7174815443338234   0.400228333963388   0.7667931773020725   0.7436575972045247   0.8219785969686663   0.453981406469929   0.29787787550642253   0.14533603116974705   0.5794543410464836   0.9727128571051609   0.6510562457440328   0.6901695263425188   0.3146405479775997   0.09727799186591488   0.22343057350377404   0.8990237911964434   0.7772431099755903   0.850491472292508   0.9907814535689815   0.2613220516752805   0.9586113972283126   0.34249556451511787   0.2689434632673539   0.45763334623966806   0.24112985289448918   0.9422672305517298   0.5021502859652813   0.7139757490351433   0.41915125592582286   0.4882858240818008   0.20427241045885883   0.5686397178653962   0.8396969148793393   0.5155729669766399   0.553216164714826   0.8784701915228775   0.5250563669017396   0.41829497511072505
0.32978559121105205   0.9794464003264342   0.7478132569261493   0.567803502818217   0.3390041376420705   0.7181243486511536   0.7892018596978367   0.22530793830309917   0.07006067437471658   0.26049100241148554   0.5480720068033476   0.28304070775136936   0.5679103884094352   0.5465152533763422   0.12892075087752464   0.7947548836695685   0.3636379779505764   0.977875535510946   0.28922383599818535   0.27918191669292863   0.8104218132357504   0.09940534398806845   0.7641674690964458   0.8608869415822036   0.4806362220246983   0.11995894366163433   0.01635421217029648   0.29308343876398657   0.14163208438262778   0.4018345950104807   0.2271523524724598   0.06777550046088737   0.0715714100079112   0.14134359259899515   0.6790803456691122   0.7847347927095181   0.503661021598476   0.5948283392226529   0.5501595947915876   0.9899799090399495   0.14002304364789958   0.6169528037117069   0.26093575879340225   0.7107979923470209   0.3296012304121493   0.5175474597236385   0.49676828969695647   0.8499110507648173   0.848965008387451   0.3975885160620042   0.48041407752666   0.5568276120008308   0.7073329240048232   0.9957539210515235   0.2532617250542002   0.4890521115399434   0.635761513996912   0.8544103284525283   0.574181379385088   0.7043173188304254   0.13210049239843602   0.2595819892298754   0.02402178459350032   0.7143374097904759
0.9920774487505365   0.6426291855181685   0.7630860258000981   0.003539417443454966   0.6624762183383872   0.12508172579452995   0.2663177361031416   0.15362836667863763   0.8135112099509362   0.7274932097325257   0.7859036585764816   0.5968007546778069   0.106178285946113   0.7317392886810022   0.5326419335222814   0.10774864313786349   0.470416771949201   0.877328960228474   0.9584605541371934   0.4034313243074381   0.338316279550765   0.6177469709985985   0.9344387695436932   0.6890939145169622   0.34623883080022855   0.97511778548043   0.1713527437435951   0.6855544970735072   0.6837626124618413   0.8500360596859001   0.9050350076404535   0.5319261303948697   0.8702514025109052   0.12254284995337437   0.11913134906397188   0.9351253757170628   0.7640731165647922   0.3908035612723721   0.5864894155416904   0.8273767325791993   0.29365634461559115   0.5134746010438982   0.628028861404497   0.42394540827176114   0.9553400650648262   0.8957276300452996   0.6935900918608038   0.7348514937547989   0.6091012342645976   0.9206098445648696   0.5222373481172087   0.04929699668129161   0.9253386218027563   0.07057378487896943   0.6172023404767552   0.5173708662864219   0.05508721929185114   0.9480309349255951   0.4980709914127833   0.5822454905693591   0.291014102727059   0.557227373653223   0.9115815758710929   0.75486875799016
0.9973577581114679   0.04375277260932481   0.28355271446659586   0.33092334971839876   0.04201769304664169   0.14802514256402519   0.5899626226057921   0.5960718559635998   0.43291645878204404   0.22741529799915564   0.0677252744885834   0.5467748592823083   0.5075778369792878   0.1568415131201862   0.45052293401182825   0.029403992995886273   0.45249061768743665   0.20881057819459115   0.952451942599045   0.44715850242652705   0.16147651496037763   0.6515832045413682   0.04087036672795208   0.6922897444363671   0.16411875684890978   0.6078304319320433   0.7573176522613562   0.3613663947179684   0.12210106380226808   0.4598052893680182   0.16735502965556412   0.7652945387543686   0.689184605020224   0.23238999136886257   0.09962975516698071   0.21851967947206033   0.18160676804093626   0.07554847824867636   0.6491068211551525   0.18911568647617405   0.7291161503534996   0.8667379000540852   0.6966548785561075   0.741957184049647   0.567639635393122   0.21515469551271704   0.6557845118281554   0.04966743961327982   0.4035208785442122   0.6073242635806737   0.8984668595667993   0.6883010448953114   0.2814198147419441   0.1475189742126555   0.7311118299112351   0.9230065061409428   0.5922352097217201   0.915128982843793   0.6314820747442544   0.7044868266688825   0.41062844168078383   0.8395805045951166   0.9823752535891019   0.5153711401927085
0.6815122913272842   0.9728426045410313   0.2857203750329944   0.7734139561430615   0.11387265593416222   0.7576879090283143   0.629935863204839   0.7237465165297817   0.71035177738995   0.15036364544764064   0.7314690036380397   0.03544547163447028   0.42893196264800587   0.0028446712349851316   0.0003571737268044642   0.11243896549352743   0.8366967529262858   0.08771568839119219   0.36887509898255   0.40795213882464487   0.426068311245502   0.2481351837960756   0.386499845393448   0.8925809986319364   0.7445560199182177   0.27529257925504425   0.10077947036045362   0.11916704248887489   0.6306833639840556   0.51760467022673   0.4708436071556147   0.3954205259590932   0.9203315865941055   0.3672410247790893   0.7393746035175751   0.3599750543246229   0.4913996239460996   0.36439635354410416   0.7390174297907706   0.24753608883109549   0.6547028710198138   0.276680665152912   0.3701423308082206   0.8395839500064506   0.22863455977431185   0.028545481356836374   0.9836424854147726   0.9470029513745142   0.4840785398560941   0.7532529021017921   0.882863015054319   0.8278359088856393   0.8533951758720386   0.23564823187506218   0.4120194078987042   0.43241538292654613   0.9330635892779331   0.8684072070959729   0.6726448043811292   0.07244032860192319   0.4416639653318335   0.5040108535518687   0.9336273745903586   0.8249042397708277
0.7869610943120197   0.22733018839895672   0.5634850437821379   0.9853202897643771   0.5583265345377079   0.19878470704212034   0.5798425583673654   0.0383173383898629   0.07424799468161374   0.44553180494032824   0.6969795433130465   0.2104814295042236   0.22085281880957516   0.20988357306526603   0.28496013541434223   0.7780660465776775   0.28778922953164204   0.34147636596929315   0.612315331033213   0.7056257179757544   0.8461252641998086   0.8374655124174245   0.6786879564428545   0.8807214782049266   0.05916416988778891   0.6101353240184677   0.11520291266071649   0.8954011884405495   0.5008376353500811   0.4113506169763474   0.535360354293351   0.8570838500506865   0.42658964066846733   0.9658188120360192   0.8383808109803046   0.646602420546463   0.2057368218588922   0.7559352389707531   0.5534206755659624   0.8685363739687855   0.9179475923272501   0.41445887300145995   0.9411053445327493   0.16291065599303123   0.07182232812744153   0.5769933605840355   0.2624173880898949   0.2821891777881046   0.012658158239652625   0.9668580365655678   0.1472144754291784   0.3867879893475551   0.5118205228895716   0.5555074195892205   0.6118541211358273   0.5297041392968685   0.08523088222110423   0.5896886075532012   0.7734733101555227   0.8831017187504056   0.879494060362212   0.8337533685824481   0.22005263458956034   0.014565344781619997
0.9615464680349619   0.41929449558098814   0.278947290056811   0.8516546887885887   0.8897241399075204   0.8423011349969526   0.01652990196691611   0.5694655110004841   0.8770659816678678   0.8754430984313848   0.8693154265377377   0.18267752165292905   0.36524545877829623   0.3199356788421644   0.25746130540191037   0.6529733823560605   0.280014576557192   0.7302470712889632   0.4839879952463877   0.7698716636056551   0.40052051619497997   0.8964937027065151   0.2639353606568273   0.755306318824035   0.438974048160018   0.47719920712552694   0.9849880706000164   0.9036516300354462   0.5492499082524976   0.6348980721285743   0.9684581686331003   0.3341861190349621   0.6721839265846299   0.7594549736971895   0.09914274209536254   0.15150859738203304   0.3069384678063336   0.4395192948550251   0.8416814366934522   0.4985352150259725   0.026923891249141633   0.7092722235660619   0.35769344144706444   0.7286635514203175   0.6264033750541617   0.8127785208595468   0.09375808079023712   0.9733572325962825   0.18742932689414366   0.33557931373401995   0.10877001019022076   0.06970560256083619   0.6381794186416461   0.7006812416054456   0.1403118415571205   0.7355194835258742   0.9659954920570162   0.9412262679082561   0.041169099461757966   0.5840108861438411   0.6590570242506826   0.501706973053231   0.19948766276830582   0.08547567111786859
0.632133133001541   0.7924347494871691   0.8417942213212414   0.3568121196975511   0.00572975794737926   0.9796562286276221   0.7480361405310042   0.3834548871012687   0.8183004310532356   0.6440769148936022   0.6392661303407835   0.3137492845404325   0.18012101241158954   0.9433956732881567   0.498954288783663   0.5782298010145583   0.21412552035457333   0.002169405379900525   0.45778518932190504   0.9942189148707173   0.5550684961038908   0.5004624323266695   0.2582975265535992   0.9087432437528487   0.9229353631023498   0.7080276828395005   0.41650330523235785   0.5519311240552975   0.9172056051549705   0.7283714542118783   0.6684671647013536   0.16847623695402886   0.09890517410173495   0.08429453931827612   0.029201034360570113   0.8547269524135964   0.9187841616901454   0.1408988660301195   0.5302467455769071   0.27649715139903797   0.7046586413355721   0.13872946065021896   0.0724615562550021   0.2822782365283207   0.14959014523168132   0.6382670283235494   0.8141640297014029   0.373534992775472   0.22665478212933152   0.930239345484049   0.39766072446904505   0.8216038687201744   0.309449176974361   0.20186789127217059   0.7291935597676915   0.6531276317661455   0.210544002872626   0.11757335195389447   0.6999925254071213   0.7984006793525492   0.2917598411824806   0.9766744859237749   0.16974577983021422   0.5219035279535112
0.5871011998469086   0.837945025273556   0.09728422357521212   0.2396252914251905   0.4375110546152272   0.19967799695000657   0.2831201938738092   0.8660902986497185   0.2108562724858957   0.26943865146595763   0.8854594694047642   0.04448642992954415   0.9014070955115348   0.06757076019378706   0.1562659096370727   0.39135879816339864   0.6908630926389087   0.9499974082398925   0.45627338422995134   0.5929581188108495   0.3991032514564281   0.9733229223161176   0.2865276043997371   0.07105459085733826   0.8120020516095195   0.13537789704256162   0.18924338082452502   0.8314292994321477   0.37449099699429234   0.935699900092555   0.9061231869507158   0.9653390007824292   0.16363472450839667   0.6662612486265974   0.020663717545951636   0.9208525708528851   0.26222762899686197   0.5986904884328104   0.864397807908879   0.5294937726894864   0.5713645363579533   0.6486930801929177   0.4081244236789276   0.9365356538786369   0.17226128490152515   0.6753701578768001   0.12159681927919046   0.8654810630212987   0.3602592332920056   0.5399922608342385   0.9323534384546655   0.03405176358915096   0.9857682362977133   0.6042923607416835   0.02623025150394966   0.06871276280672178   0.8221335117893166   0.938031112115086   0.005566533957998024   0.14786019195383676   0.5599058827924547   0.3393406236822758   0.1411687260491191   0.6183664192643503
0.9885413464345014   0.6906475434893581   0.7330443023701915   0.6818307653857134   0.8162800615329762   0.015277385612557958   0.611447483091001   0.8163497023644147   0.4560208282409706   0.47528512477831947   0.6790940446363356   0.7822979387752638   0.47025259194325736   0.8709927640366361   0.652863793132386   0.713585175968542   0.6481190801539408   0.9329616519215499   0.6472972591743879   0.5657249840147052   0.08821319736148617   0.5936210282392741   0.5061285331252688   0.9473585647503548   0.0996718509269848   0.9029734847499161   0.7730842307550773   0.26552779936464144   0.2833917893940086   0.8876960991373581   0.1616367476640763   0.44917809700022676   0.827370961153038   0.4124109743590387   0.4825427030277407   0.666880158224963   0.3571183692097806   0.5414182103224027   0.8296789098953548   0.9532949822564211   0.7089992890558398   0.6084565584008528   0.18238165072096688   0.3875699982417159   0.6207860916943536   0.014835530161578594   0.6762531175956981   0.44021143349136105   0.5211142407673688   0.11186204541166252   0.9031688868406208   0.17468363412671956   0.23772245137336026   0.2241659462743044   0.7415321391765445   0.7255055371264928   0.4103514902203223   0.8117549719152657   0.25898943614880376   0.05862537890152976   0.05323312101054169   0.2703367615928631   0.429310526253449   0.10533039664510868
0.34423383195470186   0.6618802031920104   0.2469288755324821   0.7177603984033928   0.7234477402603483   0.6470446730304318   0.570675757936784   0.2775489649120318   0.20233349949297944   0.5351826276187692   0.6675068710961632   0.10286533078531222   0.9646110481196192   0.31101668134446486   0.9259747319196188   0.37735979365881944   0.5542595578992969   0.4992617094291991   0.666985295770815   0.3187344147572897   0.5010264368887553   0.22892494783633605   0.23767476951736605   0.213404018112181   0.15679260493405334   0.5670447446443257   0.9907458939848839   0.4956436197087882   0.4333448646737051   0.920000071613894   0.4200701360480999   0.2180946547967564   0.23101136518072563   0.38481744399512474   0.7525632649519366   0.11522932401144417   0.26640031706110645   0.0738007626506599   0.8265885330323178   0.7378695303526247   0.7121407591618095   0.5745390532214608   0.15960323726150275   0.41913511559533506   0.21111432227305435   0.34561410538512477   0.9219284677441367   0.20573109748315407   0.05432171733900103   0.7785693607407991   0.9311825737592527   0.7100874777743659   0.620976852665296   0.8585692891269051   0.5111124377111529   0.4919928229776095   0.38996548748457033   0.4737518451317803   0.7585491727592163   0.3767634989661653   0.12356517042346386   0.3999510824811204   0.9319606397268985   0.6388939686135405
0.4114244112616543   0.8254120292596596   0.7723574024653957   0.2197588530182055   0.20031008898859995   0.47979792387453485   0.850428934721259   0.01402775553505142   0.1459883716495989   0.7012285631337358   0.9192463609620063   0.30394027776068555   0.525011518984303   0.8426592740068307   0.4081339232508534   0.8119474547830761   0.13504603149973263   0.36890742887505046   0.6495847504916371   0.4351839558169107   0.011480861076268773   0.96895634639393   0.7176241107647386   0.7962899872033702   0.6000564498146145   0.14354431713427046   0.9452667082993429   0.5765311341851647   0.3997463608260145   0.6637463932597356   0.0948377735780839   0.5625033786501132   0.2537579891764156   0.9625178301259998   0.17559141261607764   0.2585631008894277   0.7287464701921127   0.11985855611916901   0.7674574893652243   0.4466156461063517   0.59370043869238   0.7509511272441185   0.11787273887358712   0.011431690289440955   0.5822195776161112   0.7819947808501885   0.4002486281088485   0.2151417030860708   0.9821631278014967   0.6384504637159181   0.45498191980950553   0.6386105689009062   0.5824167669754823   0.9747040704561825   0.3601441462314216   0.07610719025079295   0.32865877779906666   0.012186240330182669   0.184552733615344   0.8175440893613652   0.599912307606954   0.8923276842110137   0.41709524425011973   0.37092844325501356
0.0062118689145739744   0.1413765569668951   0.2992225053765326   0.3594967529655726   0.4239922912984627   0.35938177611670663   0.8989738772676842   0.1443550498795018   0.441829163496966   0.7209313124007886   0.4439919574581786   0.5057444809785956   0.8594123965214837   0.7462272419446061   0.08384781122675698   0.4296372907278027   0.5307536187224171   0.7340410016144234   0.899295077611413   0.6120932013664374   0.9308413111154631   0.8417133174034098   0.48219983336129324   0.24116475811142388   0.9246294422008892   0.7003367604365147   0.18297732798476066   0.8816680051458513   0.5006371509024264   0.3409549843198081   0.2840034507170765   0.7373129552663494   0.05880798740546043   0.6200236719190195   0.8400114932588979   0.23156847428775382   0.1993955908839767   0.8737964299744133   0.7561636820321409   0.8019311835599512   0.6686419721615596   0.13975542835998989   0.8568686044207279   0.1898379821935137   0.7378006610460965   0.29804211095658006   0.37466877105943464   0.9486732240820898   0.8131712188452074   0.5977053505200653   0.19169144307467398   0.06700521893623854   0.312534067942781   0.2567503662002573   0.9076879923575975   0.3296922636698891   0.25372608053732054   0.6367266942812378   0.06767649909869962   0.09812378938213523   0.05433048965334383   0.7629302643068244   0.31151281706655876   0.2961926058221841
0.38568851749178423   0.6231748359468345   0.4546442126458308   0.10635462362867042   0.6478878564456877   0.3251327249902545   0.07997544158639623   0.15768139954658061   0.8347166376004803   0.7274273744701891   0.8882839985117222   0.09067618061034209   0.5221825696576994   0.47067700826993175   0.9805960061541248   0.760983916940453   0.26845648912037884   0.833950313988694   0.9129195070554251   0.6628601275583178   0.21412599946703503   0.07102004968186952   0.6014066899888664   0.3666675217361337   0.8284374819752508   0.44784521373503494   0.14676247734303557   0.2603128981074633   0.18054962552956308   0.12271248874478048   0.06678703575663934   0.10263149856088265   0.34583298792908274   0.3952851142745914   0.1785030372449171   0.011955317950540565   0.8236504182713833   0.9246081060046596   0.19790703109079233   0.2509714010100875   0.5551939291510045   0.09065779201596565   0.28498752403536715   0.5881112734517697   0.34106792968396943   0.019637742334096132   0.6835808340465007   0.22144375171563607   0.5126304477087186   0.5717925285990612   0.5368183567034652   0.9611308536081727   0.3320808221791555   0.4490800398542807   0.47003132094682587   0.8584993550472901   0.9862478342500728   0.0537949255796893   0.29152828370190875   0.8465440370967495   0.16259741597868946   0.12918681957502967   0.09362125261111644   0.595572636086662
0.607403486827685   0.03852902755906404   0.8086337285757492   0.00746136263489228   0.2663355571437156   0.018891285224967903   0.1250528945292485   0.7860176109192563   0.753705109434997   0.4470987566259067   0.5882345378257833   0.8248867573110834   0.42162428725584145   0.998018716771626   0.11820321687895748   0.9663874022637933   0.43537645300576866   0.9442237911919368   0.8266749331770488   0.11984336516704372   0.2727790370270792   0.815036971616907   0.7330536805659322   0.5242707290803817   0.6653755501993942   0.776507944057843   0.924419951990183   0.5168093664454894   0.39903999305567855   0.7576166588328751   0.7993670574609345   0.7307917555262332   0.6453348836206816   0.3105179022069684   0.21113251963515117   0.9059049982151498   0.22371059636484017   0.31249918543534233   0.09292930275619368   0.9395175959513564   0.7883341433590715   0.3682753942434056   0.26625436957914494   0.8196742307843128   0.5155551063319923   0.5532384226264986   0.5332006890132127   0.29540350170393104   0.8501795561325982   0.7767304785686555   0.6087807370230297   0.7785941352584417   0.4511395630769196   0.01911381973578045   0.8094136795620952   0.04780237973220843   0.805804679456238   0.708595917528812   0.5982811599269441   0.14189738151705866   0.5820940830913979   0.39609673209346974   0.5053518571707504   0.2023797855657022
0.7937599397323263   0.0278213378500641   0.2390974875916054   0.38270555478138946   0.2782048334003339   0.47458291522356555   0.7058967985783927   0.08730205307745842   0.42802527726773576   0.6978524366549099   0.09711606155536302   0.3087079178190168   0.9768857141908162   0.6787386169191295   0.2877023819932678   0.26090553808680833   0.17108103473457814   0.9701426993903175   0.6894212220663238   0.11900815656974968   0.5889869516431803   0.5740459672968478   0.18406936489557343   0.9166283710040475   0.795227011910854   0.5462246294467836   0.944971877303968   0.533922816222658   0.51702217851052   0.0716417142232181   0.23907507872557532   0.4466207631451996   0.08899690124278431   0.37378927756830815   0.1419590171702123   0.1379128453261828   0.11211118705196817   0.6950506606491786   0.8542566351769445   0.8770073072393745   0.9410301523173901   0.7249079612588611   0.1648354131106207   0.7579991506696248   0.35204320067420974   0.15086199396201344   0.9807660482150473   0.8413707796655773   0.5568161887633557   0.6046373645152298   0.03579417091107923   0.30744796344291925   0.039794010252835674   0.5329956502920117   0.7967190921855039   0.8608272002977196   0.9507971090100513   0.15920637272370358   0.6547600750152917   0.7229143549715369   0.8386859219580832   0.46415571207452494   0.8005034398383472   0.8459070477321624
0.8976557696406932   0.7392477508156639   0.6356680267277264   0.08790789706253763   0.5456125689664835   0.5883857568536504   0.6549019785126792   0.24653711739696035   0.9887963802031277   0.9837483923384206   0.6191078076015999   0.9390891539540411   0.949002369950292   0.45075274204640886   0.822388715416096   0.07826195365632144   0.9982052609402406   0.2915463693227053   0.16762864040080444   0.3553475986847846   0.15951933898215745   0.8273906572481803   0.3671252005624573   0.5094405509526222   0.2618635693414643   0.0881429064325165   0.7314571738347309   0.42153265389008454   0.7162510003749809   0.49975714957886613   0.07655519532205171   0.17499553649312422   0.7274546201718531   0.5160087572404456   0.4574473877204518   0.2359063825390831   0.7784522502215612   0.06525601519403675   0.6350586723043558   0.15764442888276167   0.7802469892813205   0.7737096458713315   0.4674300319035513   0.802296830197977   0.6207276502991631   0.9463189886231512   0.10030483134109401   0.2928562792453549   0.3588640809576988   0.8581760821906347   0.3688476575063631   0.8713236253552703   0.6426130805827179   0.3584189326117685   0.29229246218431143   0.6963280888621461   0.9151584604108647   0.8424101753713229   0.8348450744638597   0.460421706323063   0.1367062101893035   0.7771541601772862   0.1997864021595039   0.3027772774403013
0.356459220907983   0.0034445143059547026   0.7323563702559526   0.5004804472423242   0.7357315706088199   0.05712552568280353   0.6320515389148585   0.20762416799696934   0.37686748965112116   0.19894944349216886   0.26320388140849543   0.336300542641699   0.7342544090684032   0.8405305108804003   0.970911419224184   0.6399724537795529   0.8190959486575385   0.9981203355090774   0.1360663447603244   0.17955074745648986   0.682389738468235   0.22096617533179125   0.9362799426008205   0.8767734700161885   0.32593051756025204   0.21752166102583656   0.2039235723448679   0.3762930227738643   0.5901989469514322   0.16039613534303301   0.5718720334300094   0.16866885477689494   0.21333145730031097   0.9614466918508642   0.3086681520215139   0.8323683121351959   0.4790770482319077   0.12091618097046379   0.3377567327973298   0.19239585835564307   0.6599810995743692   0.12279584546138636   0.20169038803700545   0.01284511089915322   0.9775913611061342   0.9018296701295951   0.26541044543618497   0.1360716408829647   0.6516608435458822   0.6843080091037586   0.06148687309131704   0.7597786181091004   0.06146189659445   0.5239118737607256   0.4896148396613077   0.5911097633322054   0.848130439294139   0.5624651819098614   0.18094668763979385   0.7587414511970095   0.3690533910622313   0.4415490009393976   0.8431899548424641   0.5663455928413664
0.7090722914878621   0.31875315547801125   0.6414995668054586   0.5535004819422132   0.7314809303817279   0.41692348534841617   0.37608912136927364   0.41742884105924855   0.07982008683584582   0.7326154762446576   0.3146022482779566   0.6576502229501481   0.01835819024139582   0.20870360248393205   0.8249874086166489   0.06654045961794265   0.1702277509472568   0.6462384205740707   0.644040720976855   0.3077990084209331   0.8011743598850255   0.20468941963467305   0.800850766134391   0.7414534155795667   0.09210206839716344   0.8859362641566618   0.15935119932893244   0.1879529336373535   0.3606211380154355   0.46901277880824566   0.7832620779596589   0.770524092578105   0.2808010511795897   0.736397302563588   0.4686598296817022   0.11287386962795685   0.26244286093819386   0.527693700079656   0.6436724210650534   0.04633341001001421   0.09221510999093706   0.8814552795055853   0.9996317000881983   0.7385344015890811   0.2910407501059115   0.6767658598709123   0.19878093395380733   0.9970809860095143   0.1989386817087481   0.7908295957142505   0.039429734624874924   0.8091280523721609   0.8383175436933126   0.32181681690600483   0.2561676566652161   0.03860395979405594   0.5575164925137229   0.5854195143424168   0.787507826983514   0.9257300901660991   0.29507363157552907   0.057725814262760744   0.14383540591846056   0.8793966801560849
0.202858521584592   0.17627053475717536   0.1442037058302622   0.1408622785670038   0.9118177714786805   0.49950467488626304   0.9454227718764548   0.14378129255748942   0.7128790897699324   0.7086750791720126   0.90599303725158   0.3346532401853285   0.8745615460766198   0.38685826226600767   0.6498253805863639   0.2960492803912726   0.31704505356289686   0.8014387479235908   0.8623175536028499   0.3703191902251735   0.021971421987367828   0.7437129336608301   0.7184821476843893   0.4909225100690886   0.8191129004027758   0.5674423989036548   0.5742784418541271   0.3500602315020848   0.9072951289240954   0.06793772401739173   0.6288556699776723   0.20627893894459537   0.19441603915416297   0.35926264484537923   0.7228626327260924   0.8716256987592669   0.3198544930775432   0.9724043825793716   0.07303725213972855   0.5755764183679943   0.0028094395146463095   0.1709656346557807   0.21071969853687864   0.2052572281428208   0.9808380175272785   0.4272527009949506   0.49223755085248927   0.7143347180737322   0.16172511712450266   0.8598103020912958   0.9179591089983621   0.3642744865716474   0.2544299882004073   0.7918725780739041   0.2891034390206898   0.157995547627052   0.06001394904624431   0.43260993322852487   0.5662408062945975   0.28636984886778516   0.7401594559687011   0.4602055506491533   0.4932035541548689   0.7107934304997908
0.7373500164540548   0.28923991599337256   0.2824838556179903   0.50553620235697   0.7565119989267763   0.861987214998422   0.7902463047655011   0.7912014842832379   0.5947868818022737   0.0021769129071261724   0.8722871957671389   0.4269269977115905   0.3403568936018664   0.21030433483322208   0.5831837567464491   0.26893145008453845   0.2803429445556221   0.7776944016046972   0.016942950451851634   0.9825616012167533   0.540183488586921   0.3174888509555439   0.5237393962969827   0.27176817071696246   0.8028334721328662   0.028248934962171342   0.24125554067899246   0.7662319683599924   0.04632147320608982   0.16626171996374936   0.45100923591349146   0.9750304840767545   0.45153459140381613   0.16408480705662318   0.5787220401463525   0.548103486365164   0.11117769780194975   0.9537804722234011   0.9955382833999035   0.27917203628062565   0.8308347532463276   0.17608607061870388   0.9785953329480518   0.2966104350638723   0.2906512646594067   0.8585972196631599   0.4548559366510691   0.02484226434690985   0.48781779252654056   0.8303482847009886   0.21360039597207664   0.2586102959869174   0.44149631932045075   0.6640865647372393   0.7625911600585852   0.2835798119101629   0.9899617279166346   0.500001757680616   0.18386911991223265   0.7354763255449988   0.8787840301146849   0.546221285457215   0.1883308365123292   0.45630428926437316
0.04794927686835719   0.37013521483851114   0.2097355035642774   0.15969385420050086   0.7572980122089505   0.5115379951753511   0.7548795669132082   0.134851589853591   0.2694802196824099   0.6811897104743625   0.5412791709411316   0.8762412938666736   0.8279839003619592   0.017103145737123276   0.7786880108825465   0.5926614819565107   0.8380221724453246   0.5171013880565072   0.5948188909703138   0.8571851564115119   0.9592381423306398   0.9708801025992921   0.4064880544579846   0.4008808671471387   0.9112888654622826   0.600744887760781   0.1967525508937072   0.24118701294663786   0.1539908532533321   0.08920689258542992   0.4418729839804989   0.10633542309304685   0.8845106335709221   0.4080171821110674   0.9005938130393673   0.23009412922637326   0.05652673320896292   0.3909140363739441   0.12190580215682083   0.6374326472698626   0.2185045607636383   0.8738126483174369   0.5270869111865071   0.7802474908583507   0.2592664184329985   0.9029325457181447   0.12059885672852248   0.379366623711212   0.347977552970716   0.30218765795736363   0.9238463058348153   0.13817961076457413   0.1939866997173839   0.21298076537193372   0.48197332185431635   0.03184418767152729   0.3094760661464617   0.8049635832608664   0.581379508814949   0.801750058445154   0.2529493329374988   0.41404954688692225   0.45947370665812826   0.16431741117529142
0.034444772173860536   0.5402368985694853   0.9323867954716212   0.3840699203169407   0.775178353740862   0.6373043528513406   0.8117879387430987   0.004703296605728732   0.42720080077014605   0.33511669489397694   0.8879416329082834   0.8665236858411546   0.23321410105276216   0.12213592952204322   0.4059683110539671   0.8346794981696273   0.9237380349063004   0.3171723462611769   0.824588802239018   0.0329294397244733   0.6707887019688016   0.9031227993742547   0.3651150955808897   0.8686120285491818   0.636343929794941   0.36288590080476935   0.43272830010926855   0.48454210823224114   0.8611655760540791   0.7255815479534288   0.6209403613661698   0.47983881162651243   0.433964775283933   0.39046485305945183   0.7329987284578864   0.6133151257853579   0.20075067423117085   0.2683289235374086   0.32703041740391925   0.7786356276157305   0.2770126393248704   0.9511565772762317   0.5024416151649013   0.7457061878912572   0.6062239373560688   0.04803377790197708   0.13732651958401154   0.8770941593420754   0.9698800075611278   0.6851478770972077   0.704598219474743   0.3925520511098342   0.10871443150704878   0.9595663291437789   0.08365785810857321   0.9127132394833217   0.6747496562231158   0.5691014760843272   0.35065912965068685   0.29939811369796393   0.47399898199194496   0.3007725525469185   0.023628712246767585   0.5207624860822334
0.19698634266707452   0.3496159752706868   0.5211870970818663   0.7750562981909762   0.5907624053110057   0.30158219736870967   0.3838605774978548   0.8979621388489009   0.6208823977498779   0.6164343202715019   0.6792623580231117   0.5054100877390667   0.5121679662428291   0.656867991127723   0.5956044999145386   0.592696848255745   0.8374183100197133   0.08776651504339587   0.24494537026385169   0.293298734557781   0.36341932802776833   0.7869939624964774   0.2213166580170841   0.7725362484755476   0.16643298536069384   0.43737798722579063   0.7001295609352178   0.9974799502845714   0.5756705800496882   0.13579578985708096   0.31626898343736304   0.09951781143567048   0.9547881822998103   0.519361469585579   0.6370066254142512   0.5941077236966038   0.4426202160569813   0.8624934784578561   0.04140212549971273   0.001410875440858877   0.605201906037268   0.7747269634144601   0.796456755235861   0.7081121408830778   0.24178257800949965   0.9877330009179828   0.5751400972187769   0.9355758924075304   0.0753495926488058   0.5503550136921922   0.8750105362835591   0.938095942122959   0.4996790125991176   0.4145592238351112   0.5587415528461961   0.8385781306872885   0.5448908302993073   0.8951977542495322   0.9217349274319449   0.24447040699068467   0.10227061424232595   0.03270427579167616   0.8803328019322321   0.24305953154982582
0.49706870820505794   0.257977312377216   0.08387604669637105   0.5349473906667479   0.2552861301955583   0.2702443114592332   0.5087359494775942   0.5993714982592175   0.17993653754675248   0.7198892977670411   0.633725413194035   0.6612755561362587   0.6802575249476349   0.3053300739319299   0.07498386034783892   0.8226974254489702   0.13536669464832765   0.4101323196823977   0.15324893291589411   0.5782270184582855   0.03309608040600171   0.3774280438907216   0.272916130983662   0.33516748690845966   0.5360273722009438   0.11945073151350556   0.18904008428729097   0.8002200962417118   0.28074124200538547   0.8492064200542724   0.6803041348096969   0.20084859798249413   0.10080470445863297   0.12931712228723122   0.04657872161566181   0.5395730418462356   0.42054717951099807   0.8239870483553013   0.9715948612678229   0.7168756163972654   0.28518048486267045   0.41385472867290357   0.8183459283519288   0.13864859793897993   0.2520844044566687   0.036426684782182014   0.5454297973682668   0.8034811110305203   0.7160570322557249   0.9169759532686764   0.3563897130809758   0.0032610147888085497   0.43531579025033945   0.06776953321440413   0.6760855782712789   0.8024124168063144   0.3345110857917065   0.9384524109271729   0.6295068566556171   0.2628393749600789   0.9139639062807084   0.11446536257187158   0.6579119953877942   0.5459637585628135
0.628783421418038   0.7006106338989679   0.8395660670358654   0.4073151606238336   0.37669901696136926   0.664183949116786   0.29413626966759876   0.6038340495933133   0.6606419847056444   0.7472079958481095   0.937746556586623   0.6005730348045047   0.22532619445530486   0.6794384626337054   0.261660978315344   0.7981606179981904   0.8908151086635984   0.7409860517065325   0.6321541216597268   0.5353212430381115   0.9768512023828899   0.626520689134661   0.9742421262719326   0.9893574844752979   0.34806778096485197   0.9259100552356929   0.1346760592360671   0.5820423238514644   0.9713687640034827   0.26172610611890695   0.8405397895684683   0.978208274258151   0.3107267792978383   0.5145181102707974   0.9027932329818453   0.3776352394536463   0.08540058484253346   0.8350796476370921   0.6411322546665014   0.5794746214554559   0.1945854761789351   0.09409359593055956   0.008978133006774493   0.044153378417344506   0.21773427379604515   0.46757290679589864   0.03473600673484189   0.05479589394204657   0.8696664928311931   0.5416628515602057   0.9000599474987748   0.4727535700905822   0.8982977288277105   0.2799367454412987   0.059520157930306426   0.4945452958324312   0.5875709495298722   0.7654186351705012   0.15672692494846105   0.11691005637878486   0.5021703646873387   0.9303389875334092   0.5155946702819597   0.5374354349233289
0.3075848885084036   0.8362453916028496   0.5066165372751852   0.4932820565059844   0.08985061471235849   0.368672484806951   0.4718805305403433   0.4384861625639378   0.2201841218811653   0.8270096332467454   0.5718205830415685   0.9657325924733556   0.3218863930534548   0.5470728878054466   0.5123004251112621   0.47118729664092446   0.7343154435235826   0.7816542526349454   0.35557350016280104   0.3542772402621396   0.2321450788362439   0.8513152651015362   0.8399788298808414   0.8168418053388107   0.9245601903278403   0.015069873498686603   0.3333622926056562   0.3235597488328263   0.8347095756154818   0.6463973886917356   0.8614817620653129   0.8850735862688884   0.6145254537343166   0.8193877554449903   0.2896611790237444   0.9193409937955329   0.2926390606808617   0.27231486763954366   0.7773607539124823   0.4481536971546084   0.5583236171572791   0.4906606150045983   0.42178725374968123   0.09387645689246883   0.3261785383210352   0.639345349903062   0.5818084238688398   0.27703465155365814   0.4016183479931949   0.6242754764043754   0.24844613126318368   0.9534749027208318   0.5669087723777131   0.9778780877126398   0.3869643691978708   0.06840131645194336   0.9523833186433966   0.15849033226764955   0.09730319017412643   0.14906032265641048   0.6597442579625349   0.8861754646281059   0.31994243626164415   0.700906625501802
0.1014206408052558   0.39551484962350764   0.8981551825119629   0.6070301686093332   0.7752421024842207   0.7561694997204456   0.3163467586431231   0.3299955170556751   0.3736237544910257   0.13189402331607014   0.06790062737993942   0.37652061433484324   0.8067149821133126   0.1540159356034303   0.6809362581820686   0.3081192978828999   0.854331663469916   0.9955256033357808   0.5836330680079422   0.1590589752264894   0.1945874055073811   0.10935013870767488   0.26369063174629803   0.4581523497246873   0.0931667647021253   0.7138352890841673   0.3655354492343351   0.8511221811153541   0.3179246622179047   0.9576657893637217   0.049188690591211996   0.521126664059679   0.944300907726879   0.8257717660476516   0.9812880632112726   0.14460604972483576   0.13758592561356642   0.6717558304442213   0.30035180502920394   0.8364867518419359   0.2832542621436504   0.6762302271084405   0.7167187370212618   0.6774277766154465   0.08866685663626932   0.5668800884007655   0.45302810527496373   0.21927542689075916   0.995500091934144   0.8530447993165984   0.08749265604062861   0.36815324577540504   0.6775754297162393   0.8953790099528767   0.03830396544941662   0.8470265817157261   0.7332745219893603   0.06960724390522514   0.05701590223814404   0.7024205319908903   0.5956885963757939   0.39785141346100394   0.7566640972089401   0.8659337801489544
0.31243433423214345   0.7216211863525634   0.03994536018767835   0.18850600353350788   0.22376747759587415   0.15474109795179788   0.5869172549127146   0.9692305766427487   0.22826738566173013   0.30169629863519953   0.499424598872086   0.6010773308673436   0.5506919559454908   0.40631728868232286   0.4611206334226694   0.7540507491516176   0.8174174339561305   0.3367100447770977   0.4041047311845254   0.05163021716072736   0.22172883758033662   0.9388586313160938   0.6474406339755853   0.185696437011773   0.9092945033481932   0.2172374449635303   0.6074952737879069   0.9971904334782651   0.685527025752319   0.06249634701173245   0.02057801887519228   0.027959856835516397   0.4572596400905889   0.7608000483765329   0.5211534200031063   0.4268825259681727   0.906567684145098   0.35448275969421006   0.06003278658043682   0.6728317768165551   0.08915025018896754   0.017772714917112346   0.6559280553959115   0.6212015596558278   0.8674214126086309   0.07891408360101856   0.008487421420326161   0.4355051226440548   0.9581269092604378   0.8616766386374882   0.40099214763241925   0.43831468916578964   0.2725998835081187   0.7991802916257558   0.38041412875722697   0.41035483233027326   0.8153402434175299   0.03838024324922288   0.8592607087541208   0.9834723063621005   0.9087725592724317   0.6838974835550128   0.7992279221736839   0.3106405295455454
0.8196223090834642   0.6661247686379005   0.14329986677777246   0.6894389698897176   0.9522008964748333   0.5872106850368819   0.1348124453574463   0.25393384724566287   0.9940739872143955   0.7255340463993937   0.7338202977250271   0.8156191580798733   0.7214741037062768   0.9263537547736379   0.3534061689678001   0.4052643257496   0.906133860288747   0.8879735115244151   0.4941454602136794   0.4217920193874995   0.9973613010163153   0.2040760279694022   0.6949175380399955   0.11115148984195407   0.177738991932851   0.5379512593315017   0.551617671262223   0.4217125199522364   0.2255380954580177   0.9507405742946198   0.41680522590477675   0.16777867270657354   0.23146410824362212   0.2252065278952261   0.6829849281797498   0.3521595146267003   0.5099900045373452   0.2988527731215882   0.3295787592119496   0.9468951888771003   0.6038561442485982   0.4108792615971732   0.8354332989982702   0.5251031694896009   0.606494843232283   0.20680323362777103   0.14051576095827473   0.4139516796476468   0.428755851299432   0.6688519742962693   0.5888980896960517   0.9922391596954103   0.2032177558414143   0.7181114000016495   0.17209286379127492   0.8244604869888368   0.9717536475977921   0.4929048721064234   0.4891079356115252   0.4723009723621365   0.4617636430604469   0.19405209898483516   0.1595291763995756   0.5254057834850362
0.8579074988118487   0.783172837387662   0.32409587740130535   0.0003026139954353175   0.25141265557956566   0.5763696037598909   0.18358011644303063   0.5863509343477885   0.8226568042801337   0.9075176294636216   0.5946820267469789   0.5941117746523782   0.6194390484387193   0.1894062294619721   0.42258916295570403   0.7696512876635414   0.6476854008409272   0.6965013573555487   0.9334812273441788   0.2973503153014049   0.1859217577804803   0.5024492583707135   0.7739520509446032   0.7719445318163687   0.3280142589686317   0.7192764209830516   0.4498561735432978   0.7716419178209334   0.076601603389066   0.14290681722316065   0.2662760571002672   0.18529098347314485   0.25394479910893236   0.23538918775953901   0.6715940303532882   0.5911792088207667   0.634505750670213   0.04598295829756692   0.24900486739758426   0.8215279211572253   0.9868203498292858   0.3494816009420182   0.3155236400534055   0.5241776058558204   0.8008985920488054   0.8470323425713047   0.5415715891088023   0.7522330740394517   0.4728843330801738   0.1277559215882531   0.09171541556550444   0.9805911562185183   0.3962827296911078   0.9848491043650924   0.8254393584652372   0.7953001727453735   0.14233793058217545   0.7494599166055534   0.15384532811194898   0.20412096392460682   0.5078321799119625   0.7034769583079865   0.9048404607143647   0.38259304276738154
0.5210118300826767   0.3539953573659683   0.5893168206609593   0.8584154369115611   0.7201132380338713   0.5069630147946637   0.047745231552156965   0.10618236287210939   0.2472289049536975   0.3792070932064105   0.9560298159866525   0.12559120665359105   0.8509461752625898   0.39435798884131806   0.13059045752141527   0.33029103390821757   0.7086082446804143   0.6448980722357647   0.9767451294094663   0.12617006998361072   0.20077606476845183   0.941421113927778   0.0719046686951016   0.7435770272162292   0.6797642346857751   0.5874257565618098   0.48258784803414234   0.8851615903046681   0.9596509966519038   0.08046274176714618   0.4348426164819854   0.7789792274325587   0.7124220916982063   0.7012556485607356   0.47881280049533287   0.6533880207789676   0.8614759164356165   0.3068976597194176   0.34822234297391763   0.32309698687075006   0.15286767175520222   0.661999587483653   0.3714772135644513   0.19692691688713937   0.9520916069867504   0.7205784735558749   0.2995725448693497   0.45334988967091017   0.2723273723009753   0.13315271699406508   0.8169846968352074   0.5681882993662422   0.3126763756490715   0.05268997522691891   0.38214208035322195   0.7892090719336834   0.6002542839508652   0.35143432666618324   0.903329279857889   0.1358210511547158   0.7387783675152487   0.04453666694676562   0.5551069368839714   0.8127240642839657
0.5859106957600465   0.3825370794631126   0.18362972331952016   0.6157971473968263   0.6338190887732961   0.6619586059072378   0.8840571784501704   0.1624472577259162   0.3614917164723208   0.5288058889131726   0.06707248161496313   0.5942589583596741   0.048815340823249266   0.4761159136862537   0.6849304012617412   0.8050498864259906   0.448561056872384   0.1246815870200705   0.7816011214038522   0.6692288352712749   0.7097826893571353   0.08014492007330488   0.2264941845198807   0.8565047709873091   0.12387199359708875   0.6976078406101922   0.042864461200360554   0.24070762359048276   0.49005290482379266   0.03564923470295453   0.1588072827501901   0.07826036586456656   0.12856118835147184   0.5068433457897819   0.09173480113522699   0.48400140750489246   0.07974584752822259   0.03072743210352815   0.4068043998734858   0.6789515210789018   0.6311847906558385   0.9060458450834576   0.6252032784696336   0.009722685807626964   0.9214021012987033   0.8259009250101528   0.39870909394975296   0.15321791482031785   0.7975301077016146   0.1282930843999605   0.3558446327493924   0.9125102912298351   0.3074772028778219   0.09264384969700598   0.1970373499992023   0.8342499253652685   0.17891601452635006   0.585800503907224   0.1053025488639753   0.3502485178603761   0.09917016699812746   0.5550730718036959   0.6984981489904895   0.6712969967814743
0.4679853763422889   0.6490272267202383   0.07329487052085584   0.6615743109738473   0.5465832750435856   0.8231263017100855   0.6745857765711029   0.5083563961535295   0.749053167341971   0.694833217310125   0.3187411438217105   0.5958461049236944   0.44157596446414915   0.602189367613119   0.1217037938225082   0.7615961795584258   0.2626599499377991   0.016388863705894933   0.016401244958532894   0.41134766169804976   0.16348978293967162   0.461315791902199   0.3179030959680434   0.7400506649165756   0.6955044065973828   0.8122885651819607   0.24460822544718755   0.07847635394272823   0.14892113155379716   0.9891622634718752   0.5700224488760847   0.5701199577891988   0.39986796421182613   0.29432904616175015   0.2512813050543742   0.9742738528655044   0.958291999747677   0.6921396785486311   0.12957751123186595   0.21267767330707862   0.6956320498098779   0.6757508148427361   0.11317626627333306   0.8013300116090288   0.5321422668702063   0.2144350229405372   0.7952731703052897   0.061279346692453336   0.8366378602728235   0.4021464577585765   0.5506649448581021   0.9828029927497252   0.6877167287190263   0.41298419428670136   0.9806424959820175   0.41268303496052633   0.28784876450720026   0.11865514812495119   0.7293611909276433   0.4384091820950219   0.3295567647595233   0.4265154695763201   0.5997836796957774   0.22573150878794326
0.6339247149496454   0.7507646547335839   0.4866074134224443   0.4244014971789144   0.10178244807943918   0.5363296317930467   0.6913342431171546   0.36312215048646107   0.2651445878066157   0.13418317403447017   0.14066929825905247   0.38031915773673597   0.5774278590875893   0.7211989797477688   0.160026802277035   0.9676361227762097   0.2895790945803891   0.6025438316228177   0.4306656113493917   0.5292269406811878   0.9600223298208659   0.17602836204649755   0.8308819316536143   0.3034954318932445   0.3260976148712204   0.4252637073129137   0.34427451823117006   0.8790939347143301   0.22431516679178123   0.888934075519867   0.6529402751140154   0.515971784227869   0.9591705789851656   0.7547509014853968   0.5122709768549629   0.13565262649113302   0.3817427198975762   0.033551921737628   0.35224417457792795   0.16801650371492335   0.0921636253171871   0.4310080901148104   0.9215785632285363   0.6387895630337356   0.13214129549632125   0.2549797280683128   0.09069663157492193   0.33529413114049106   0.8060436806251008   0.8297160207553992   0.7464221133437519   0.45620019642616094   0.5817285138333196   0.9407819452355322   0.09348183822973642   0.9402284121982919   0.622557934848154   0.18603104375013535   0.5812108613747735   0.8045757857071589   0.2408152149505778   0.15247912201250735   0.2289666867968455   0.6365592819922355
0.14865158963339073   0.721471031897697   0.30738812356830925   0.9977697189585   0.016510294137069458   0.46649130382938414   0.2166914919933873   0.6624755878180089   0.21046661351196863   0.636775283073985   0.4702693786496354   0.20627539139184795   0.628738099678649   0.6959933378384529   0.376787540419899   0.266046979193556   0.006180164830495025   0.5099622940883175   0.7955766790451255   0.4614711934863971   0.7653649498799172   0.3574831720758101   0.56660999224828   0.8249119114941615   0.6167133602465265   0.6360121401781131   0.2592218686799708   0.8271421925356616   0.6002030661094571   0.16952083634872897   0.04253037668658352   0.16466660471765265   0.3897364525974884   0.5327455532747439   0.5722609980369481   0.9583912133258047   0.7609983529188393   0.8367522154362911   0.1954734576170491   0.6923442341322487   0.7548181880883443   0.32678992134797363   0.3998967785719235   0.2308730406458516   0.9894532382084271   0.9693067492721635   0.8332867863236435   0.4059611291516901   0.3727398779619006   0.3332946090940504   0.5740649176436726   0.5788189366160285   0.7725368118524436   0.16377377274532143   0.5315345409570892   0.4141523318983758   0.3828003592549552   0.6310282194705775   0.959273542920141   0.4557611185725711   0.6218020063361158   0.7942760040342863   0.763800085303092   0.7634168844403224
0.8669838182477715   0.4674860826863127   0.36390330673116844   0.5325438437944708   0.8775305800393444   0.49817933341414916   0.5306165204075249   0.12658271464278076   0.5047907020774437   0.16488472432009874   0.9565516027638523   0.5477637780267522   0.7322538902250002   0.001110951574777307   0.4250170618067632   0.13361144612837644   0.349453530970045   0.37008273210419984   0.46574351888662213   0.6778503275558053   0.7276515246339291   0.5758067280699135   0.7019434335835302   0.9144334431154829   0.8606677063861576   0.1083206453836008   0.33804012685236173   0.38188959932101213   0.9831371263468133   0.6101413119694516   0.8074236064448368   0.25530688467823137   0.4783464242693696   0.4452565876493529   0.8508720036809845   0.7075431066514791   0.7460925340443694   0.4441456360745756   0.42585494187422135   0.5739316605231026   0.3966390030743244   0.07406290397037577   0.9601114229875992   0.8960813329672973   0.6689874784403953   0.4982561759004623   0.25816798940406904   0.9816478898518144   0.8083197720542376   0.3899355305168615   0.9201278625517073   0.5997582905308023   0.8251826457074243   0.7797942185474098   0.11270425610687052   0.34445140585257095   0.34683622143805476   0.33453763089805694   0.26183225242588604   0.6369082992010918   0.6007436873936853   0.8903919948234813   0.8359773105516647   0.06297663867798918
0.20410468431936094   0.8163290908531056   0.8758658875640655   0.16689530571069183   0.5351172058789657   0.3180729149526433   0.6176978981599964   0.1852474158588774   0.7267974338247281   0.9281373844357819   0.6975700356082891   0.5854891253280751   0.9016147881173038   0.148343165888372   0.5848657795014186   0.24103771947550415   0.5547785666792491   0.813805534990315   0.32303352707553257   0.6041294202744123   0.9540348792855637   0.9234135401668337   0.4870562165238679   0.5411527815964231   0.7499301949662027   0.10708444931372815   0.6111903289598024   0.37425747588573127   0.21481298908723706   0.7890115343610848   0.993492430799806   0.18901006002685386   0.488015555262509   0.860874149925303   0.29592239519151686   0.6035209346987788   0.5864007671452052   0.712530984036931   0.7110566156900983   0.3624832152232746   0.03162220046595613   0.898725449046616   0.3880230886145657   0.7583537949488623   0.07758732118039244   0.9753119088797823   0.9009668720906978   0.21720101335243922   0.3276571262141897   0.8682274595660541   0.2897765431308954   0.8429435374667079   0.11284413712695261   0.07921592520496924   0.2962841123310894   0.6539334774398541   0.6248285818644437   0.21834177527966622   0.0003617171395725162   0.05041254274107532   0.038427814719238444   0.5058107912427352   0.28930510144947424   0.6879293275178007
0.006805614253282315   0.6070853421961192   0.9012820128349085   0.9295755325689384   0.9292182930728898   0.631773433316337   0.0003151407442107039   0.7123745192164992   0.6015611668587002   0.7635459737502829   0.7105385976133153   0.8694309817497913   0.4887170297317476   0.6843300485453137   0.4142544852822259   0.21549750430993717   0.863888447867304   0.46598827326564746   0.4138927681426534   0.16508496156886185   0.8254606331480655   0.9601774820229123   0.12458766669317917   0.47715563405106115   0.8186550188947832   0.35309213982679305   0.22330565385827064   0.5475801014821228   0.8894367258218934   0.721318706510456   0.22299051311405993   0.8352055822656236   0.2878755589631931   0.9577727327601732   0.5124519155007446   0.9657746005158323   0.7991585292314455   0.2734426842148595   0.09819743021851872   0.7502770962058952   0.9352700813641416   0.8074544109492121   0.6843046620758654   0.5851921346370333   0.10980944821607605   0.8472769289262998   0.5597169953826862   0.1080365005859722   0.2911544293212928   0.49418478909950675   0.33641134152441554   0.5604563991038495   0.4017177034993995   0.7728660825890507   0.11342082841035558   0.7252508168382259   0.11384214453620639   0.8150933498288775   0.600968912909611   0.7594762163223935   0.31468361530476086   0.541650665614018   0.5027714826910923   0.009199120116498356
0.37941353394061933   0.734196254664806   0.8184668206152269   0.424006985479465   0.26960408572454325   0.8869193257385062   0.25874982523254075   0.31597048489349283   0.9784496564032504   0.3927345366389994   0.9223384837081252   0.7555140857896434   0.5767319529038509   0.6198684540499487   0.8089176552977696   0.030263268951417545   0.4628898083676445   0.8047751042210711   0.20794874238815866   0.270787052629024   0.14820619306288363   0.26312443860705315   0.7051772596970665   0.26158793251252566   0.7687926591222644   0.5289281839422472   0.8867104390818396   0.8375809470330606   0.49918857339772105   0.642008858203741   0.6279606138492988   0.5216104621395677   0.5207389169944706   0.2492743215647416   0.7056221301411736   0.7660963763499243   0.9440069640906197   0.6294058675147929   0.896704474843404   0.7358331073985068   0.4811171557229752   0.8246307632937218   0.6887557324552452   0.46504605476948285   0.33291096266009157   0.5615063246866686   0.9835784727581788   0.20345812225695717   0.5641183035378272   0.03257814074442142   0.0968680336763393   0.3658771752238965   0.0649297301401062   0.3905692825406804   0.4689074198270405   0.8442667130843288   0.5441908131456356   0.1412949609759388   0.763285289685867   0.07817033673440435   0.6001838490550159   0.5118890934611459   0.866580814842463   0.3423372293358975
0.1190666933320406   0.6872583301674242   0.17782508238721775   0.8772911745664147   0.786155730671949   0.12575200548075557   0.19424660962903892   0.6738330523094576   0.22203742713412178   0.09317386473633414   0.09737857595269962   0.307955877085561   0.15710769699401558   0.7026045821956537   0.6284711561256591   0.4636891640012322   0.6129168838483801   0.561309621219715   0.8651858664397921   0.3855188272668279   0.012733034793364191   0.04942052775856903   0.9986050515973292   0.04318159793093037   0.8936663414613236   0.3621621975911449   0.8207799692101114   0.1658904233645157   0.10751061078937456   0.2364101921103893   0.6265333595810725   0.4920573710550582   0.8854731836552527   0.14323632737405514   0.5291547836283729   0.1841014939694972   0.7283654866612372   0.4406317451784014   0.9006836275027138   0.720412329968265   0.11544860281285718   0.8793221239586865   0.035497761062921615   0.33489350270143714   0.102715568019493   0.8299015962001175   0.036892709465592456   0.29171190477050674   0.2090492265581694   0.46773939860897257   0.21611274025548105   0.12582148140599106   0.10153861576879486   0.2313292064985833   0.5895793806744085   0.6337641103509328   0.21606543211354207   0.08809287912452814   0.06042459704603565   0.4496626163814357   0.4876999454523049   0.6474611339461267   0.15974096954332187   0.7292502864131707
0.3722513426394477   0.7681390099874402   0.12424320848040026   0.39435678371173355   0.2695357746199547   0.9382374137873227   0.08735049901480779   0.1026448789412268   0.06048654806178527   0.47049801517835016   0.8712377587593267   0.9768233975352357   0.9589479322929905   0.2391688086797669   0.2816583780849182   0.3430592871843029   0.7428825001794483   0.15107592955523877   0.22123378103888258   0.8933966708028672   0.25518255472714346   0.503614795609112   0.06149281149556071   0.16414638438969656   0.8829312120876958   0.7354757856216718   0.9372496030151605   0.769789600677963   0.6133954374677411   0.7972383718343491   0.8498991040003526   0.6671447217367362   0.5529088894059558   0.3267403566559989   0.9786613452410259   0.6903213242015005   0.5939609571129654   0.08757154797623197   0.6970029671561077   0.3472620370171976   0.851078456933517   0.9364956184209932   0.4757691861172251   0.4538653662143304   0.5958959022063736   0.43288082281188117   0.4142763746216644   0.28971898182463385   0.7129646901186778   0.6974050371902093   0.4770267716065039   0.5199293811466708   0.09956925265093669   0.9001666653558603   0.6271276676061512   0.8527846594099345   0.5466603632449809   0.5734263086998614   0.6484663223651254   0.1624633352084341   0.9526994061320154   0.48585476072362943   0.9514633552090177   0.8152012981912364
0.10162094919849837   0.5493591423026363   0.47569416909179263   0.3613359319769061   0.5057250469921248   0.11647831949075507   0.06141779447012823   0.07161695015227228   0.792760356873447   0.41907328230054575   0.5843910228636243   0.5516875690056015   0.6931911042225103   0.5189066169446854   0.9572633552574731   0.6989029095956669   0.14653074097752944   0.945480308244824   0.3087970328923477   0.5364395743872328   0.19383133484551401   0.4596255475211946   0.35733367768333   0.7212382761959963   0.09221038564701563   0.9102664052185584   0.8816395085915374   0.3599023442190902   0.5864853386548908   0.7937880857278033   0.8202217141214092   0.2882853940668179   0.7937249817814438   0.3747148034272576   0.23583069125778486   0.7365978250612164   0.10053387755893353   0.8558081864825722   0.2785673360003118   0.03769491546554957   0.9540031365814041   0.9103278782377481   0.9697703031079641   0.5012553410783168   0.76017180173589   0.45070233071655347   0.6124366254246341   0.7800170648823205   0.6679614160888745   0.5404359254979951   0.7307971168330967   0.4201147206632303   0.0814760774339836   0.7466478397701918   0.9105754027116876   0.1318293265964124   0.28775109565253976   0.37193303634293423   0.6747447114539027   0.39523150153519593   0.18721721809360622   0.5161248498603621   0.3961773754535909   0.35753658606964633
0.23321408151220213   0.605796971622614   0.4264070723456268   0.8562812449913295   0.4730422797763121   0.1550946409060605   0.8139704469209927   0.07626418010900908   0.8050808636874376   0.6146587154080654   0.083173330087896   0.6561494594457787   0.723604786253454   0.8680108756378736   0.17259792737620847   0.5243201328493664   0.4358536906009142   0.49607783929493937   0.4978532159223058   0.12908863131417048   0.248636472507308   0.9799529894345773   0.1016758404687149   0.7715520452445241   0.015422390995105874   0.37415601781196334   0.6752687681230881   0.9152708002531945   0.5423801112187938   0.2190613769059028   0.8612983212020954   0.8390066201441855   0.7372992475313562   0.6044026614978374   0.7781249911141994   0.18285716069840668   0.013694461277902217   0.7363917858599638   0.6055270637379909   0.6585370278490403   0.577840770676988   0.24031394656502444   0.10767384781568513   0.5294483965348699   0.32920429816968   0.26036095713044716   0.005998007346970228   0.7578963512903457   0.3137819071745741   0.8862049393184839   0.3307292392238821   0.8426255510371512   0.7714017959557803   0.667143562412581   0.4694309180217867   0.003618930892965675   0.03410254842442407   0.0627409009147436   0.6913059269075873   0.820761770194559   0.020408087146521852   0.32634911505477976   0.08577886316959635   0.16222474234551867
0.44256731646953384   0.08603516848975536   0.9781050153539113   0.6327763458106489   0.1133630182998539   0.8256742113593082   0.9721070080069409   0.8748799945203032   0.7995811111252799   0.9394692720408244   0.6413777687830589   0.032254443483152005   0.028179315169499522   0.2723257096282434   0.17194685076127217   0.02863551259018633   0.9940767667450755   0.2095848087134998   0.4806409238536849   0.20787374239562736   0.9736686795985536   0.88323569365872   0.3948620606840885   0.04564900005010867   0.5311013631290197   0.7972005251689647   0.4167570453301773   0.4128726542394598   0.41773834482916583   0.9715263138096564   0.4446500373232363   0.5379926597191567   0.618157233703886   0.03205704176883203   0.8032722685401774   0.5057382162360047   0.5899779185343865   0.7597313321405886   0.6313254177789053   0.4771027036458183   0.595901151789311   0.5501465234270888   0.1506844939252204   0.26922896125019097   0.6222324721907575   0.6669108297683689   0.7558224332411319   0.2235799612000823   0.09113110906173773   0.8697103045994042   0.33906538791095453   0.8107073069606224   0.6733927642325719   0.8981839907897478   0.8944153505877181   0.2727146472414658   0.055235530528685864   0.8661269490209158   0.09114308204754071   0.7669764310054612   0.4652576119942993   0.10639561688032712   0.4598176642686354   0.28987372735964284
0.8693564602049882   0.5562490934532383   0.30913317034341503   0.02064476610945188   0.24712398801423083   0.8893382636848695   0.5533107371022832   0.7970648049093696   0.1559928789524931   0.0196279590854652   0.21424534919132865   0.986357497948747   0.4826001147199212   0.12144396829571742   0.31982999860361044   0.7136428507072813   0.42736458419123535   0.25531701927480166   0.22868691655606976   0.9466664197018201   0.962106972196936   0.14892140239447457   0.7688692522874343   0.6567926923421772   0.09275051199194771   0.5926723089412363   0.4597360819440193   0.6361479262327253   0.8456265239777169   0.7033340452563669   0.9064253448417361   0.8390831213233557   0.6896336450252237   0.6837060861709017   0.6921799956504074   0.8527256233746087   0.20703353030530255   0.5622621178751843   0.372349997046797   0.1390827726673274   0.7796689461140672   0.3069450986003826   0.14366308049072726   0.19241635296550733   0.8175619739171313   0.15802369620590803   0.37479382820329293   0.5356236606233301   0.7248114619251835   0.5653513872646717   0.9150577462592736   0.8994757343906047   0.8791849379474667   0.8620173420083048   0.008632401417537463   0.06039261306724896   0.18955129292224288   0.17831125583740315   0.31645240576712996   0.20766698969264027   0.9825177626169403   0.6160491379622188   0.9441024087203329   0.06858421702531287
0.2028488165028731   0.3091040393618363   0.8004393282296057   0.8761678640598055   0.38528684258574186   0.15108034315592825   0.42564550002631274   0.34054420343647546   0.6604753806605583   0.5857289558912565   0.5105877537670391   0.4410684690458707   0.7812904427130917   0.7237116138829517   0.5019553523495017   0.38067585597862175   0.5917391497908489   0.5454003580455485   0.18550294658237174   0.1730088662859815   0.6092213871739085   0.9293512200833296   0.24140053786203877   0.10442464926066862   0.40637257067103544   0.6202471807214933   0.44096120963243307   0.22825678520086307   0.021085728085293576   0.4691668375655651   0.015315709606120338   0.8877125817643876   0.36061034742473524   0.8834378816743086   0.5047279558390811   0.4466441127185169   0.5793199047116435   0.15972626779135693   0.0027726034895794944   0.06596825673989513   0.9875807549207947   0.6143259097458084   0.8172696569072078   0.8929593904539136   0.3783593677468862   0.6849746896624788   0.575869119045169   0.7885347411932451   0.9719867970758508   0.0647275089409854   0.1349079094127359   0.560277955992382   0.9509010689905572   0.5955606713754203   0.11959219980661556   0.6725653742279943   0.590290721565822   0.7121227897011118   0.6148642439675344   0.22592126150947742   0.010970816854178408   0.5523965219097547   0.6120916404779548   0.1599530047695823
0.023390061933383693   0.9380706121639464   0.7948219835707471   0.26699361431566865   0.6450306941864975   0.2530959225014676   0.2189528645255781   0.47845887312242363   0.6730438971106467   0.1883684135604822   0.08404495511284221   0.9181809171300417   0.7221428281200896   0.5928077421850619   0.9644527553062267   0.24561554290204737   0.1318521065542676   0.8806849524839502   0.3495885113386923   0.019694281392569936   0.12088128970008918   0.32828843057419543   0.7374968708607375   0.8597412766229876   0.09749122776670549   0.39021781841024905   0.9426748872899903   0.592747662307319   0.452460533580208   0.1371218959087814   0.7237220227644122   0.11428878918489534   0.7794166364695613   0.9487534823482991   0.63967706765157   0.19610787205485367   0.057273808349471725   0.35594574016323727   0.6752243123453433   0.9504923291528062   0.9254217017952041   0.4752607876792871   0.325635801006651   0.9307980477602363   0.804540412095115   0.14697235710509168   0.5881389301459136   0.07105677113724872   0.7070491843284095   0.7567545386948427   0.6454640428559233   0.4783091088299297   0.2545886507482015   0.6196326427860612   0.9217420200915112   0.3640203196450344   0.4751720142786402   0.670879160437762   0.2820649524399412   0.16791244759018073   0.4178982059291685   0.3149334202745247   0.6068406400945978   0.21742011843737444
0.4924765041339643   0.8396726325952376   0.28120483908794686   0.2866220706771381   0.6879360920388494   0.692700275490146   0.6930659089420332   0.2155652995398894   0.98088690771044   0.9359457367953034   0.04760186608610992   0.7372561907099596   0.7262982569622385   0.3163130940092421   0.1258598459945988   0.3732358710649253   0.2511262426835983   0.64543393357148   0.8437948935546576   0.20532342347474453   0.8332280367544298   0.3305005132969554   0.23695425346005974   0.9879033050373701   0.3407515326204655   0.49082788070171773   0.9557494143721129   0.7012812343602319   0.6528154405816161   0.7981276052115718   0.2626835054300796   0.4857159348203426   0.6719285328711762   0.8621818684162684   0.21508163934396973   0.748459744110383   0.9456302759089377   0.5458687744070263   0.08922179334937094   0.3752238730454577   0.6945040332253394   0.9004348408355463   0.24542689979471333   0.16990044957071315   0.8612759964709096   0.5699343275385909   0.008472646334653602   0.1819971445333431   0.520524463850444   0.07910644683687314   0.052723231962540716   0.4807159101731111   0.8677090232688279   0.28097884162530135   0.790039726532461   0.9949999753527685   0.19578049039765177   0.4187969732090329   0.5749580871884914   0.24654023124238558   0.25015021448871405   0.8729281988020066   0.4857362938391204   0.8713163581969279
0.5556461812633746   0.9724933579664603   0.24030939404440707   0.7014159086262147   0.694370184792465   0.4025590304278694   0.23183674770975346   0.5194187640928717   0.17384572094202097   0.32345258359099627   0.17911351574721274   0.038702853919760576   0.306136697673193   0.04247374196569492   0.38907378921475166   0.043702878566992044   0.11035620727554125   0.623676768756662   0.8141157020262604   0.7971626473246064   0.8602059927868272   0.7507485699546554   0.3283794081871399   0.9258462891276785   0.3045598115234526   0.7782552119881951   0.08807001414273286   0.22443038050146374   0.6101896267309875   0.37569618156032575   0.8562332664329794   0.7050116164085921   0.43634390578896654   0.05224359796932948   0.6771197506857667   0.6663087624888315   0.13020720811577352   0.00976985600363456   0.28804596147101497   0.6226058839218395   0.019851000840232252   0.38609308724697255   0.47393025944475464   0.825443236597233   0.15964500805340506   0.6353445172923171   0.14555085125761474   0.8995969474695544   0.8550851965299525   0.8570893053041219   0.057480837114881875   0.6751665669680907   0.24489556979896498   0.48139312374379617   0.20124757068190247   0.9701549505594986   0.8085516640099984   0.4291495257744667   0.5241278199961358   0.30384618807066716   0.678344455894225   0.41937966977083213   0.23608185852512084   0.6812403041488277
0.6584934550539927   0.03328658252385956   0.7621515990803662   0.8557970675515947   0.4988484470005876   0.39794206523154246   0.6166007478227514   0.9562001200820403   0.6437632504706352   0.5408527599274205   0.5591199107078696   0.2810335531139495   0.39886768067167017   0.059459636183624445   0.35787234002596713   0.3108786025544508   0.5903160166616718   0.6303101104091577   0.8337445200298312   0.007032414483783679   0.9119715607674468   0.21093044063832567   0.5976626615047105   0.325792110334956   0.2534781057134541   0.17764385811446612   0.8355110624243443   0.4699950427833613   0.7546296587128665   0.7797017928829236   0.21891031460159277   0.5137949227013211   0.1108664082422313   0.23884903295550303   0.6597904038937232   0.2327613695873716   0.7119987275705612   0.1793893967718786   0.3019180638677561   0.9218827670329207   0.12168271090888941   0.5490792863627209   0.4681735438379248   0.914850352549137   0.20971115014144262   0.33814884572439513   0.8705108823332144   0.5890582422141811   0.9562330444279885   0.16050498760992904   0.0349998199088701   0.11906319943081982   0.20160338571512207   0.3808031947270054   0.8160895053072773   0.6052682767294988   0.09073697747289078   0.14195416177150239   0.15629910141355413   0.37250690714212714   0.3787382499023296   0.9625647649996237   0.8543810375457981   0.4506241401092064
0.25705553899344025   0.413485478636903   0.3862074937078733   0.5357737875600693   0.047344388851997626   0.07533663291250783   0.5156966113746589   0.9467155453458882   0.09111134442400909   0.9148316453025788   0.4806967914657888   0.8276523459150684   0.889507958708887   0.5340284505755734   0.6646072861585115   0.22238406918556963   0.7987709812359962   0.392074288804071   0.5083081847449574   0.8498771620434425   0.4200327313336666   0.42950952380444724   0.6539271471991593   0.3992530219342361   0.16297719234022634   0.016024045167544257   0.26771965349128607   0.8634792343741668   0.11563280348822873   0.9406874122550364   0.7520230421166272   0.9167636890282786   0.024521459064219632   0.02585576695245761   0.2713262506508384   0.08911134311321028   0.1350135003553326   0.4918273163768842   0.6067189644923269   0.8667272739276406   0.3362425191193364   0.0997530275728132   0.09841077974736948   0.016850111884198153   0.9162097877856697   0.670243503768366   0.44448363254821016   0.617597089949962   0.7532325954454434   0.6542194586008216   0.17676397905692406   0.7541178555757952   0.6375997919572147   0.7135320463457853   0.4247409369402969   0.8373541665475166   0.6130783328929951   0.6876762793933276   0.15341468628945854   0.7482428234343063   0.47806483253766247   0.19584896301644344   0.5466957217971317   0.8815155495066657
0.14182231341832607   0.09609593544363026   0.4482849420497622   0.8646654376224675   0.2256125256326563   0.4258524316752643   0.0038013095015520916   0.24706834767250543   0.47237993018721286   0.7716329730744427   0.827037330444628   0.4929504920967102   0.8347801382299982   0.05810092672865735   0.40229639350433116   0.6555963255491937   0.22170180533700312   0.3704246473353297   0.2488817072148726   0.9073535021148874   0.7436369727993407   0.17457568431888623   0.7021859854177409   0.025837952608221797   0.6018146593810145   0.07847974887525597   0.2539010433679787   0.16117251498575433   0.37620213374835826   0.6526273171999917   0.2500997338664266   0.914104167313249   0.9038222035611454   0.880994344125549   0.42306240342179857   0.4211536752165387   0.0690420653311472   0.8228934173968917   0.020766009917467406   0.765557349667345   0.8473402599941441   0.452468770061562   0.7718843027025948   0.8582038475524576   0.10370328719480343   0.2778930857426758   0.06969831728485391   0.8323658949442357   0.5018886278137888   0.1994133368674198   0.8157972739168753   0.6711933799584814   0.1256864940654306   0.5467860196674281   0.5656975400504487   0.7570892126452325   0.22186429050428522   0.6657916755418791   0.14263513662865013   0.33593553742869386   0.152822225173138   0.8428982581449874   0.12186912671118272   0.5703781877613489
0.3054819651789939   0.3904294880834254   0.3499848240085879   0.7121743402088914   0.2017786779841905   0.11253640234074963   0.280286506723734   0.8798084452646555   0.6998900501704016   0.9131230654733298   0.4644892328068587   0.20861506530617413   0.574203556104971   0.3663370458059017   0.89879169275641   0.4515258526609416   0.35233926560068585   0.7005453702640225   0.75615655612776   0.11559031523224772   0.1995170404275478   0.8576471121190351   0.6342874294165772   0.5452121274708989   0.8940350752485539   0.46721762403560974   0.28430260540798935   0.8330377872620075   0.6922563972643634   0.3546812216948601   0.0040160986842553365   0.953229341997352   0.9923663470939618   0.4415581562215303   0.5395268658773966   0.7446142766911777   0.41816279098899073   0.07522111041562861   0.6407351731209865   0.2930884240302362   0.06582352538830492   0.37467574015160604   0.8845786169932266   0.17749810879798847   0.8663064849607571   0.5170286280325709   0.2502911875766493   0.6322859813270897   0.9722714097122033   0.049811003996961124   0.96598858216866   0.7992481940650822   0.28001501244783983   0.695129782302101   0.9619724834844047   0.8460188520677302   0.28764866535387806   0.2535716260805707   0.4224456176070081   0.10140457537655241   0.8694858743648873   0.1783505156649421   0.7817104444860216   0.8083161513463162
0.8036623489765824   0.8036747755133361   0.897131827492795   0.6308180425483277   0.9373558640158253   0.28664614748076517   0.6468406399161457   0.998532061221238   0.965084454303622   0.23683514348380405   0.6808520577474857   0.19928386715615595   0.6850694418557822   0.5417053611817031   0.718879574263081   0.3532650150884257   0.3974207765019042   0.2881337351011323   0.29643395665607286   0.25186043971187333   0.5279349021370169   0.10978321943619024   0.5147235121700513   0.4435442883655571   0.7242725531604345   0.3061084439228542   0.6175916846772563   0.8127262458172294   0.7869166891446092   0.019462296442089008   0.9707510447611106   0.8141941845959912   0.8218322348409872   0.782627152958285   0.28989898701362504   0.6149103174398354   0.136762792985205   0.24092179177658193   0.571019412750544   0.2616453023514096   0.7393420164833008   0.9527880566754496   0.27458545609447116   0.009784862639536283   0.2114071143462839   0.8430048372392593   0.7598619439244199   0.5662405742739792   0.48713456118584936   0.5368963933164052   0.14227025924716352   0.7535143284567498   0.7002178720412401   0.5174340968743162   0.17151921448605284   0.9393201438607586   0.8783856372002529   0.7348069439160312   0.8816202274724279   0.32440982642092325   0.7416228442150479   0.4938851521394493   0.3106008147218837   0.06276452406951366
0.0022808277317470896   0.5410970954639996   0.036015358627412564   0.05297966142997737   0.7908737133854632   0.6980922582247403   0.2761534147029927   0.4867390871559982   0.30373915219961384   0.16119586490833518   0.1338831554558292   0.7332247586992483   0.6035212801583737   0.643761768034019   0.9623639409697764   0.7939046148384897   0.7251356429581208   0.9089548241179878   0.08074371349734856   0.46949478841756653   0.983512798743073   0.41506967197853856   0.7701428987754648   0.4067302643480529   0.9812319710113259   0.8739725765145389   0.7341275401480523   0.35375060291807553   0.19035825762586267   0.1758803182897985   0.45797412544505955   0.8670115157620774   0.8866191054262489   0.014684453381463342   0.3240909699892303   0.13378675706282897   0.28309782526787514   0.3709226853474443   0.36172702901945397   0.3398821422243392   0.5579621823097543   0.46196786122945654   0.2809833155221054   0.8703873538067727   0.5744493835666813   0.046898189250917995   0.5108404167466406   0.4636570894587198   0.5932174125553554   0.17292561273637916   0.7767128765985883   0.10990648654064428   0.4028591549294928   0.9970452944465806   0.3187387511535288   0.24289497077856695   0.516240049503244   0.9823608410651173   0.9946477811642984   0.10910821371573799   0.23314222423536884   0.611438155717673   0.6329207521448444   0.7692260714913988
0.6751800419256145   0.14947029448821644   0.3519374366227391   0.8988387176846262   0.1007306583589332   0.10257210523729844   0.8410970198760985   0.43518162822590634   0.5075132458035777   0.9296464925009192   0.06438414327751017   0.32527514168526206   0.10465409087408492   0.9326011980543386   0.7456453921239814   0.08238017090669512   0.588414041370841   0.9502403569892214   0.7509976109596829   0.9732719571909572   0.3552718171354721   0.3388022012715484   0.11807685881483841   0.20404588569955834   0.6800917752098575   0.18933190678333198   0.7661394221920993   0.3052071680149322   0.5793611168509244   0.08675980154603352   0.9250424023160008   0.8700255397890259   0.07184787104734665   0.15711330904511422   0.8606582590384906   0.5447503981037638   0.9671937801732617   0.22451211099077556   0.11501286691450925   0.4623702271970686   0.3787797388024208   0.27427175400155424   0.36401525595482637   0.4890982700061115   0.023507921666948664   0.9354695527300058   0.2459383971399879   0.28505238430655316   0.34341614645709106   0.7461376459466739   0.4797989749478886   0.9798452162916209   0.7640550296061667   0.6593778444006403   0.5547565726318878   0.10981967650259512   0.6922071585588201   0.5022645353555261   0.6940983135933971   0.5650692783988314   0.7250133783855583   0.2777524243647505   0.579085446678888   0.10269905120176276
0.3462336395831375   0.0034806703631963163   0.21507019072406156   0.6136007811956513   0.32272571791618887   0.06801111763319051   0.9691317935840736   0.32854839688909815   0.9793095714590978   0.32187347168651664   0.48933281863618505   0.3487031805974772   0.21525454185293108   0.6624956272858763   0.9345762460042972   0.23888350409488204   0.523047383294111   0.16023109193035026   0.2404779324109001   0.6738142256960507   0.7980340049085527   0.8824786675655998   0.6613924857320121   0.571115174494288   0.4518003653254152   0.8789979972024035   0.4463222950079506   0.9575143932986366   0.1290746474092263   0.8109868795692129   0.477190501423877   0.6289659964095385   0.14976507595012853   0.48911340788269625   0.9878576827876919   0.2802628158120613   0.9345105340971974   0.8266177805968199   0.053281436783394726   0.041379311717179276   0.41146315080308643   0.6663866886664697   0.8128035043724946   0.36756508602112864   0.6134291458945338   0.7839080211008699   0.15141101864048245   0.7964499115268407   0.16162878056911856   0.9049100238984665   0.7050887236325318   0.8389355182282041   0.03255413315989226   0.0939231443292536   0.22789822220865483   0.2099695218186656   0.8827890572097638   0.6048097364465573   0.24004053942096287   0.9297067060066043   0.9482785231125663   0.7781919558497374   0.18675910263756815   0.888327394289425
0.5368153723094798   0.11180526718326783   0.3739555982650735   0.5207623082682964   0.923386226414946   0.3278972460823979   0.22254457962459104   0.7243123967414556   0.7617574458458275   0.4229872221839314   0.5174558559920592   0.8853768785132515   0.7292033126859353   0.32906407785467784   0.2895576337834044   0.675407356694586   0.8464142554761716   0.7242543414081205   0.0495170943624415   0.7457006506879816   0.8981357323636052   0.9460623855583831   0.8627579917248733   0.8573732563985567   0.36132036005412543   0.8342571183751152   0.48880239345979987   0.33661094813026027   0.4379341336391793   0.5063598722927173   0.2662578138352088   0.6122985513888045   0.6761766877933518   0.08337265010878585   0.7488019578431496   0.726921672875553   0.9469733751074165   0.754308572254108   0.45924432405974525   0.051514316180967024   0.10055911963124493   0.030054230845987535   0.40972722969730374   0.30581366549298533   0.20242338726763967   0.08399184528760452   0.5469692379724304   0.4484404090944287   0.8411030272135143   0.24973472691248932   0.05816684451263054   0.11182946096416845   0.4031688935743349   0.743374854619772   0.7919090306774217   0.4995309095753639   0.7269922057809831   0.6600022045109862   0.04310707283427211   0.7726092366998109   0.7800188306735667   0.9056936322568782   0.5838627487745268   0.7210949205188438
0.6794597110423217   0.8756394014108907   0.1741355190772231   0.4152812550258585   0.477036323774682   0.7916475561232862   0.6271662811047928   0.9668408459314298   0.6359332965611678   0.5419128292107969   0.5689994365921622   0.8550113849672614   0.2327644029868329   0.7985379745910247   0.7770904059147404   0.3554804753918975   0.5057721972058498   0.13853577008003856   0.7339833330804684   0.5828712386920866   0.7257533665322832   0.23284213782316038   0.1501205843059415   0.8617763181732427   0.046293655489961415   0.35720273641226974   0.9759850652287184   0.4464950631473842   0.5692573317152794   0.5655551802889835   0.34881878412392564   0.47965421721595436   0.9333240351541116   0.02364235107818676   0.7798193475317634   0.624642832248693   0.7005596321672787   0.225104376487162   0.002728941617023   0.2691623568567955   0.19478743496142886   0.08656860640712344   0.26874560853655466   0.686291118164709   0.46903406842914575   0.8537264685839631   0.11862502423061316   0.8245147999914663   0.4227404129391843   0.4965237321716933   0.1426399590018948   0.378019736844082   0.8534830812239049   0.9309685518827098   0.7938211748779691   0.8983655196281276   0.9201590460697934   0.907326200804523   0.014001827346205696   0.2737226873794346   0.21959941390251475   0.682221824317361   0.011272885729182695   0.0045603305226391
0.0248119789410859   0.5956532179102376   0.742527277192628   0.31826921235793015   0.5557779105119401   0.7419267493262746   0.6239022529620148   0.4937544123664639   0.13303749757275585   0.24540301715458115   0.4812622939601201   0.11573467552238188   0.2795544163488509   0.3144344652718714   0.6874411190821509   0.21736915589425423   0.3593953702790575   0.4071082644673484   0.6734392917359452   0.9436464685148196   0.13979595637654274   0.7248864401499874   0.6621664060067626   0.9390861379921804   0.11498397743545685   0.1292332222397498   0.9196391288141345   0.6208169256342503   0.5592060669235167   0.3873064729134753   0.2957368758521196   0.12706251326778642   0.4261685693507608   0.14190345575889413   0.8144745818919995   0.011327837745404544   0.1466141530019099   0.8274689904870227   0.1270334628098486   0.7939586818511504   0.7872187827228524   0.42036072601967434   0.4535941710739034   0.8503122133363308   0.6474228263463097   0.695474285869687   0.7914277650671409   0.9112260753441502   0.5324388489108528   0.5662410636299372   0.8717886362530064   0.2904091497098999   0.9732327819873361   0.17893459071646187   0.5760517604008868   0.16334663644211347   0.5470642126365753   0.03703113495756774   0.7615771785088872   0.15201879869670895   0.4004500596346654   0.209562144470545   0.6345437156990387   0.3580601168455586
0.613231276911813   0.7892014184508707   0.18094954462513524   0.5077479035092279   0.9658084505655034   0.09372713258118369   0.3895217795579944   0.5965218281650776   0.4333696016546505   0.5274860689512465   0.5177331433049881   0.30611267845517776   0.4601368196673144   0.34855147823478466   0.9416813829041013   0.14276604201306425   0.9130726070307391   0.3115203432772169   0.18010420439521407   0.9907472433163553   0.5126225473960737   0.1019581988066719   0.5455604886961755   0.6326871264707967   0.8993912704842607   0.31275678035580123   0.3646109440710402   0.12493922296156879   0.9335828199187574   0.21902964777461756   0.9750891645130458   0.5284173947964912   0.5002132182641068   0.691543578823371   0.4573560212080578   0.2223047163413134   0.04007639859679247   0.34299210058858637   0.5156746383039564   0.07953867432824915   0.1270037915660534   0.031471757311369475   0.3355704339087424   0.08879143101189385   0.6143812441699797   0.9295135585046975   0.790009945212567   0.4561043045410972   0.714989973685719   0.6167567781488963   0.4253990011415267   0.3311650815795284   0.7814071537669617   0.39772713037427876   0.4503098366284809   0.8027476867830372   0.2811939355028549   0.7061835515509077   0.992953815420423   0.5804429704417239   0.24111753690606239   0.36319145096232136   0.4772791771164666   0.5009042961134746
0.11411374534000898   0.3317196936509519   0.14170874320772422   0.41211286510158085   0.49973250117002926   0.4022061351462543   0.3516987979951573   0.9560085605604837   0.7847425274843102   0.785449356997358   0.9262997968536306   0.6248434789809553   0.0033353737173484766   0.3877222266230792   0.4759899602251497   0.8220957921979181   0.7221414382144936   0.6815386750721715   0.4830361448047266   0.2416528217561942   0.4810239013084312   0.31834722410985006   0.00575696768826001   0.7407485256427195   0.36691015596842225   0.9866275304588982   0.8640482244805358   0.3286356605411387   0.867177654798393   0.5844213953126438   0.5123494264853785   0.372627099980655   0.08243512731408281   0.7989720383152858   0.5860496296317479   0.7477836209996997   0.07909975359673432   0.41124981169220665   0.1100596694065982   0.9256878288017817   0.3569583153822407   0.7297111366200352   0.6270235246018716   0.6840350070455875   0.8759344140738095   0.4113639125101851   0.6212665569136115   0.943286481402868   0.5090242581053873   0.42473638205128694   0.7572183324330758   0.6146508208617293   0.6418466033069943   0.8403149867386431   0.24486890594769728   0.24202372088107424   0.5594114759929115   0.041342948423357256   0.6588192763159494   0.49424009988137446   0.48031172239617714   0.6300931367311506   0.5487596069093511   0.5685522710795927
0.12335340701393642   0.9003820001111155   0.9217360823074796   0.8845172640340052   0.24741899294012693   0.4890180876009303   0.300469525393868   0.9412307826311372   0.7383947348347397   0.06428170554964337   0.5432511929607922   0.3265799617694079   0.0965481315277454   0.22396671881100025   0.29838228701309494   0.08455624088833368   0.5371366555348339   0.182623770387643   0.6395630106971456   0.5903161410069592   0.05682493313865679   0.5525306336564924   0.09080340378779445   0.02176386992736645   0.9334715261247204   0.652148633545377   0.16906732148031486   0.13724660589336124   0.6860525331845935   0.16313054594444665   0.8685977960864469   0.19601582326222403   0.9476577983498538   0.09884884039480328   0.32534660312565467   0.869435861492816   0.8511096668221084   0.8748821215838031   0.02696431611255973   0.7848796206044825   0.31397301128727445   0.6922583511961601   0.3874013054154141   0.19456347959752324   0.2571480781486177   0.13972771753966765   0.2965979016276197   0.17279960967015678   0.3236765520238973   0.4875790839942907   0.12753058014730484   0.035553003776795544   0.6376240188393039   0.324448538049844   0.25893278406085796   0.8395371805145715   0.6899662204894501   0.22559969765504076   0.9335861809352033   0.9701013190217554   0.8388565536673417   0.3507175760712377   0.9066218648226435   0.185221698417273
0.5248835423800673   0.6584592248750777   0.5192205594072294   0.9906582188197498   0.2677354642314496   0.5187315073354101   0.22262265777960968   0.817858609149593   0.9440589122075523   0.031152423341119374   0.09509207763230487   0.7823056053727975   0.3064348933682484   0.7067038852912754   0.8361592935714469   0.942768424858226   0.6164686728787984   0.4811041876362346   0.9025731126362436   0.9726671058364705   0.7776121192114566   0.13038661156499684   0.9959512478136001   0.7874454074191974   0.25272857683138933   0.4719273866899191   0.47673068840637073   0.7967871885994477   0.9849931125999397   0.9531958793545091   0.254108030626761   0.9789285794498547   0.04093420039238743   0.9220434560133897   0.15901595299445614   0.1966229740770572   0.734499307024139   0.21533957072211438   0.32285665942300923   0.25385454921883127   0.11803063414534068   0.7342353830858798   0.42028354678676555   0.2811874433823608   0.3404185149338841   0.603848771520883   0.42433229897316543   0.4937420359631633   0.08768993810249474   0.13192138483096383   0.9476016105667947   0.6969548473637156   0.10269682550255502   0.17872550547645474   0.6934935799400337   0.7180262679138609   0.061762625110167585   0.25668204946306505   0.5344776269455775   0.5214032938368037   0.3272633180860286   0.041342478740950685   0.21162096752256834   0.26754874461797246
0.20923268394068792   0.3071070956550709   0.7913374207358027   0.9863613012356116   0.8688141690068039   0.703258324134188   0.3670051217626373   0.49261926527244837   0.781124230904309   0.5713369393032242   0.41940351119584257   0.7956644179087328   0.6784274054017541   0.39261143382676933   0.7259099312558088   0.07763814999487188   0.6166647802915864   0.1359293843637043   0.19143230431023128   0.5562348561580682   0.2894014622055579   0.09458690562275361   0.979811336787663   0.28868611154009577   0.08016877826486998   0.7874798099676827   0.1884739160518602   0.3023248103044841   0.21135460925806615   0.0842214858334948   0.8214687942892229   0.8097055450320357   0.43023037835375705   0.5128845465302707   0.40206528309338035   0.01404112712330292   0.751802972952003   0.12027311270350133   0.6761553518375715   0.936402977128431   0.13513819266041652   0.984343728339797   0.4847230475273402   0.38016812097036284   0.8457367304548586   0.8897568227170434   0.5049117107396772   0.09148200943026709   0.7655679521899886   0.10227701274936069   0.316437794687817   0.789157199125783   0.5542133429319225   0.018055526915865892   0.49496900039859415   0.9794516540937472   0.12398296457816542   0.5051709803855952   0.09290371730521381   0.9654105269704444   0.37217999162616244   0.3848978676820939   0.4167483654676423   0.029007549842013324
0.2370417989657459   0.40055413934229683   0.9320253179403021   0.6488394288716505   0.39130506851088726   0.5107973166252534   0.42711360720062486   0.5573574194413834   0.6257371163208987   0.4085203038758928   0.11067581251280782   0.7682002203156004   0.07152377338897616   0.39046477696002685   0.6157068121142136   0.7887485662218531   0.9475408088108107   0.8852937965744316   0.5228030948089999   0.8233380392514087   0.5753608171846483   0.5003959288923377   0.10605472934135755   0.7943304894093954   0.3383190182189024   0.09984178955004092   0.17402941140105543   0.14549106053774494   0.9470139497080151   0.5890444729247875   0.7469158042004306   0.5881336410963616   0.3212768333871165   0.18052416904889473   0.6362399916876228   0.8199334207807611   0.24975305999814035   0.7900593920888679   0.020533179573409083   0.031184854558908067   0.3022122511873296   0.9047655955144362   0.4977300847644092   0.20784681530749932   0.7268514340026813   0.40436966662209844   0.39167535542305165   0.4135163258981039   0.3885324157837789   0.30452787707205753   0.21764594402199622   0.268025265360359   0.4415184660757637   0.7154834041472701   0.47073013982156564   0.6798916242639974   0.12024163268864722   0.5349592350983753   0.8344901481339428   0.8599582034832363   0.8704885726905068   0.7448998430095074   0.8139569685605338   0.8287733489243282
0.5682763215031773   0.8401342474950713   0.31622688379612457   0.6209265336168288   0.8414248875004959   0.43576458087297276   0.924551528373073   0.20741020771872493   0.4528924717167171   0.13123670380091523   0.7069055843510768   0.939384942358366   0.011374005640953378   0.4157532996536452   0.23617544452951109   0.2594933180943686   0.8911323729523062   0.8807940645552699   0.4016852963955682   0.39953511461113234   0.020643800261799267   0.13589422154576242   0.5877283278350345   0.5707617656868041   0.452367478758622   0.2957599740506912   0.27150144403890986   0.9498352320699753   0.610942591258126   0.8599953931777184   0.34694991566583694   0.7424250243512504   0.1580501195414089   0.7287586893768031   0.6400443313147602   0.8030400819928845   0.1466761139004555   0.31300538972315795   0.4038688867852491   0.5435467638985159   0.25554374094814936   0.43221132516788807   0.0021835903896809013   0.1440116492873835   0.23489994068635012   0.2963171036221257   0.4144552625546465   0.5732498836005794   0.7825324619277281   0.0005571295714345021   0.14295381851573663   0.623414651530604   0.1715898706696021   0.1405617363937161   0.7960039028498997   0.8809896271793536   0.013539751128193198   0.41180304701691295   0.1559595715351395   0.07794954518646922   0.8668636372277376   0.09879765729375498   0.7520906847498904   0.5344027812879534
0.6113198962795883   0.6665863321258668   0.7499070943602095   0.3903911320005699   0.3764199555932382   0.37026922850374117   0.335451831805563   0.8171412483999906   0.5938874936655101   0.36971209893230667   0.19249801328982638   0.19372659686938654   0.42229762299590795   0.22915036253859059   0.39649411043992666   0.3127369696900329   0.4087578718677148   0.8173473155216776   0.24053453890478718   0.23478742450356369   0.5418942346399771   0.7185496582279227   0.48844385415489683   0.7003846432156103   0.9305743383603888   0.0519633261020558   0.7385367597946874   0.30999351121504043   0.5541543827671506   0.6816940975983146   0.4030849279891243   0.49285226281504985   0.9602668891016405   0.3119819986660079   0.21058691469929797   0.2991256659456633   0.5379692661057326   0.08283163612741733   0.8140928042593712   0.9863886962556304   0.12921139423801778   0.2654843206057397   0.5735582653545841   0.7516012717520667   0.5873171595980407   0.546934662377817   0.08511441119968728   0.051216628536456435   0.6567428212376519   0.49497133627576123   0.34657765140499996   0.741223117321416   0.10258843847050127   0.8132772386774466   0.9434927234158756   0.24837085450636615   0.14232154936886074   0.5012952400114387   0.7329058087165776   0.9492451885607028   0.6043522832631282   0.4184636038840214   0.9188130044572064   0.9628564923050724
0.47514088902511037   0.15297928327828167   0.3452547391026223   0.21125522055300563   0.8878237294270697   0.6060446209004646   0.260140327902935   0.1600385920165492   0.23108090818941784   0.11107328462470345   0.9135626764979351   0.4188154746951332   0.12849246971891656   0.29779604594725684   0.9700699530820595   0.17044462018876705   0.9861709203500558   0.7965008059358182   0.23716414436548175   0.22119943162806424   0.38181863708692765   0.3780372020517968   0.31835113990827535   0.25834293932299185   0.9066777480618172   0.22505791877351516   0.9730964008056531   0.04708771876998622   0.018854018634747532   0.6190132978730505   0.712956072902718   0.8870491267534371   0.7877731104453297   0.507940013248347   0.799393396404783   0.4682336520583038   0.6592806407264131   0.2101439673010902   0.8293234433227236   0.29778903186953676   0.6731097203763573   0.413643161365272   0.5921592989572418   0.0765896002414725   0.29129108328942965   0.035605959313475204   0.27380815904896644   0.8182466609184806   0.38461333522761243   0.81054804053996   0.30071175824331337   0.7711589421484945   0.3657593165928649   0.19153474266690954   0.5877556853405953   0.8841098153950574   0.5779862061475352   0.6835947294185625   0.7883622889358124   0.4158761633367536   0.918705565421122   0.4734507621174723   0.9590388456130888   0.11808713146721685
0.24559584504476473   0.05980760075220024   0.366879546655847   0.04149753122574434   0.9543047617553351   0.02420164143872504   0.09307138760688052   0.2232508703072637   0.5696914265277226   0.213653600898765   0.7923596293635672   0.45209192815876925   0.20393210993485775   0.022118858231855457   0.2046039440229718   0.5679821127637119   0.6259459037873225   0.33852412881329297   0.4162416550871595   0.15210594942695826   0.7072403383662005   0.8650733666958207   0.4572028094740707   0.03401881795974142   0.46164449332143576   0.8052657659436204   0.09032326281822373   0.9925212867339971   0.5073397315661007   0.7810641245048954   0.9972518752113432   0.7692704164267334   0.937648305038378   0.5674105236061304   0.20489224584777604   0.31717848826796413   0.7337161951035203   0.545291665374275   0.00028830182480424   0.7491963755042522   0.10777029131619777   0.20676753656098198   0.5840466467376447   0.597090426077294   0.40052995294999727   0.34169416986516127   0.12684383726357407   0.5630716081175525   0.9388854596285615   0.5364284039215408   0.036520574445350354   0.5705503213835554   0.4315457280624609   0.7553642794166454   0.039268699234007165   0.8012799049568221   0.49389742302408285   0.187953755810515   0.8343764533862311   0.484101416688858   0.7601812279205625   0.64266209043624   0.8340881515614269   0.7349050411846058
0.6524109366043648   0.43589455387525805   0.2500415048237821   0.13781461510731174   0.25188098365436745   0.09420038401009677   0.12319766756020803   0.5747430069897592   0.31299552402580594   0.5577719800885559   0.08667709311485766   0.004192685606203685   0.881449795963345   0.8024077006719105   0.047408393880850504   0.2029127806493816   0.3875523729392622   0.6144539448613955   0.2130319404946194   0.7188113639605236   0.6273711450186997   0.9717918544251555   0.3789437889331925   0.9839063227759179   0.974960208414335   0.5358973005498975   0.12890228410941043   0.8460917076686062   0.7230792247599674   0.4416969165398007   0.005704616549202398   0.271348700678847   0.41008370073416156   0.8839249364512447   0.9190275234343447   0.2671560150726433   0.5286339047708165   0.08151723577933422   0.8716191295534942   0.0642432344232617   0.14108153183155428   0.4670632909179387   0.6585871890588748   0.3454318704627381   0.5137103868128545   0.4952714364927832   0.2796434001256823   0.3615255476868202   0.5387501783985196   0.9593741359428858   0.15074111601627188   0.515433840018214   0.8156709536385521   0.5176772194030851   0.14503649946706948   0.24408513933936707   0.40558725290439057   0.6337522829518404   0.22600897603272477   0.9769291242667237   0.8769533481335741   0.5522350471725062   0.35438984647923055   0.9126858898434621
0.7358718163020198   0.08517175625456745   0.6958026574203557   0.567254019380724   0.22216142948916523   0.5899003197617843   0.4161592572946734   0.2057284716939038   0.6834112510906456   0.6305261838188985   0.2654181412784015   0.6902946316756897   0.8677402974520935   0.11284896441581341   0.12038164181133201   0.4462094923363227   0.4621530445477029   0.47909668146397305   0.8943726657786073   0.4692803680695989   0.5851996964141288   0.926861634291467   0.5399828192993767   0.5565944782261368   0.849327880112109   0.8416898780368994   0.844180161879021   0.9893404588454128   0.6271664506229438   0.25178955827511523   0.4280209045843476   0.783611987151509   0.9437551995322983   0.6212633744562167   0.1626027633059461   0.09331735547581926   0.07601490208020475   0.5084144100404033   0.042221121494614114   0.6471078631394966   0.6138618575325019   0.02931772857643024   0.14784845571600685   0.17782749506989776   0.028662161118373043   0.10245609428496331   0.6078656364166302   0.621233016843761   0.179334281006264   0.26076621624806384   0.7636854745376092   0.6318925579983482   0.5521678303833202   0.008976657972948627   0.33566456995326155   0.8482805708468392   0.6084126308510219   0.3877132835167319   0.1730618066473154   0.75496321537102   0.5323977287708171   0.8792988734763286   0.13084068515270128   0.10785535223152329
0.9185358712383154   0.8499811448998984   0.9829922294366944   0.9300278571616255   0.8898737101199423   0.747525050614935   0.3751265930200643   0.3087948403178646   0.7105394291136783   0.48675883436687123   0.6114411184824551   0.6769022823195164   0.1583715987303581   0.47778217639392256   0.2757765485291936   0.8286217114726773   0.5499589678793362   0.09006889287719066   0.1027147418818782   0.07365849610165734   0.017561239108518943   0.21077001940086207   0.9718740567291769   0.965803143870134   0.0990253678702036   0.3607888745009637   0.9888818272924825   0.0357752867085085   0.20915165775026132   0.6132638238860286   0.6137552342724182   0.726980446390644   0.49861222863658305   0.12650498951915745   0.0023141157899630727   0.0500781640711275   0.34024062990622495   0.6487228131252348   0.7265375672607695   0.22145645259845026   0.7902816620268888   0.5586539202480442   0.6238228253788912   0.14779795649679292   0.7727204229183698   0.3478839008471821   0.6519487686497144   0.1819948126266589   0.6736950550481662   0.9870950263462185   0.6630669413572319   0.14621952591815038   0.4645433972979049   0.3738312024601898   0.049311707084813694   0.4192390795275065   0.9659311686613219   0.24732621294103235   0.04699759129485062   0.36916091545637897   0.625690538755097   0.5986033998157975   0.32046002403408114   0.1477044628579287
0.8354088767282082   0.039949479567753264   0.6966371986551899   0.9999065063611358   0.0626884538098383   0.6920655787205711   0.04468843000547551   0.8179116937344769   0.38899339876167205   0.7049705523743527   0.38162148864824363   0.6716921678163265   0.9244500014637672   0.3311393499141629   0.33230978156342994   0.25245308828882   0.9585188328024453   0.08381313697313053   0.2853121902685793   0.8832921728324411   0.33282829404734837   0.48520973715733307   0.9648521662344981   0.7355877099745124   0.4974194173191402   0.44526025758957977   0.26821496757930824   0.7356812036133765   0.4347309635093019   0.7531946788690087   0.22352653757383276   0.9177695098788997   0.045737564747629834   0.04822412649465601   0.8419050489255892   0.2460773420625732   0.12128756328386267   0.7170847765804931   0.5095952673621592   0.9936242537737532   0.16276873048141738   0.6332716396073627   0.22428307709357992   0.11033208094131212   0.829940436434069   0.14806190245002954   0.25943091085908176   0.37474437096679974   0.3325210191149288   0.7028016448604497   0.9912159432797735   0.6390631673534232   0.897790055605627   0.9496069659914411   0.7676894057059408   0.7212936574745235   0.8520524908579971   0.9013828394967851   0.9257843567803516   0.4752163154119503   0.7307649275741345   0.18429806291629194   0.4161890894181924   0.4815920616381971
0.5679961970927171   0.5510264233089294   0.19190601232461246   0.37125998069688504   0.738055760658648   0.4029645208588998   0.9324751014655307   0.9965156097300852   0.40553474154371916   0.7001628759984501   0.9412591581857571   0.35745244237666207   0.5077446859380922   0.7505559100070089   0.1735697524798164   0.6361587849021385   0.6556921950800951   0.8491730705102238   0.24778539569946478   0.16094246949018826   0.9249272675059607   0.6648750075939319   0.8315963062812723   0.6793504078519911   0.3569310704132437   0.11384858428500261   0.63969029395666   0.3080904271551061   0.6188753097545957   0.7108840634261028   0.7072151924911293   0.31157481742502086   0.2133405682108765   0.010721187427652793   0.7659560343053721   0.9541223750483588   0.7055958822727842   0.2601652774206438   0.5923862818255557   0.3179635901462203   0.04990368719268915   0.41099220691041993   0.3446008861260909   0.157021120656032   0.12497641968672846   0.746117199316488   0.5130045798448185   0.4776707128040409   0.7680453492734848   0.6322686150314853   0.8733142858881585   0.1695802856489348   0.14917003951888913   0.9213845516053826   0.1660990933970293   0.8580054682239139   0.9358294713080126   0.9106633641777298   0.4001430590916572   0.9038830931755552   0.23023358903522834   0.650498086757086   0.8077567772661015   0.5859195030293348
0.1803299018425392   0.239505879846666   0.4631558911400106   0.42889838237330286   0.05535348215581074   0.493388680530178   0.950151311295192   0.951227669569262   0.28730813288232593   0.8611200654986926   0.07683702540703352   0.7816473839203272   0.13813809336343683   0.93973551389331   0.9107379320100042   0.9236419156964133   0.20230862205542421   0.02907214971558021   0.510594872918347   0.01975882252085813   0.9720750330201958   0.3785740629584943   0.7028380956522455   0.43383931949152327   0.7917451311776567   0.13906818311182828   0.2396822045122349   0.004940937118220396   0.736391649021846   0.6456795025816503   0.2895308932170428   0.05371326754895842   0.44908351613951997   0.7845594370829577   0.2126938678100093   0.27206588362863127   0.31094542277608317   0.8448239231896477   0.30195593580000507   0.34842396793221797   0.10863680072065895   0.8157517734740676   0.7913610628816581   0.3286651454113598   0.1365617677004631   0.43717771051557325   0.08852296722941257   0.8948258259198366   0.3448166365228064   0.29810952740374497   0.8488407627171777   0.8898848888016162   0.6084249875009605   0.6524300248220947   0.5593098695001348   0.8361716212526578   0.15934147136144053   0.867870587739137   0.3466160016901256   0.5641057376240265   0.8483960485853573   0.023046664549489157   0.04466006589012051   0.21568176969180855
0.7397592478646984   0.20729489107542162   0.2532990030084624   0.8870166242804487   0.6031974801642354   0.7701171805598483   0.1647760357790499   0.9921907983606121   0.2583808436414289   0.4720076531561034   0.3159352730618722   0.1023059095589959   0.6499558561404684   0.8195776283340087   0.7566254035617374   0.2661342883063381   0.49061438477902786   0.9517070405948718   0.4100094018716118   0.7020285506823116   0.6422183361936705   0.9286603760453827   0.3653493359814913   0.48634678099050305   0.902459088328972   0.721365484969961   0.11205033297302883   0.5993301567100544   0.29926160816473674   0.9512483044101127   0.9472742971939789   0.6071393583494422   0.040880764523307814   0.47924065125400933   0.6313390241321067   0.5048334487904463   0.3909249083828394   0.6596630229200006   0.8747136205703694   0.23869916048410822   0.9003105236038116   0.7079559823251288   0.4647042186987576   0.5366706098017966   0.25809218741014106   0.7792956062797461   0.09935488271726632   0.050323828811293554   0.35563309908116897   0.057930121309785136   0.9873045497442375   0.4509936721012392   0.05637149091643227   0.10668181689967246   0.04003025255025856   0.843854313751797   0.015490726393124456   0.6274411656456631   0.4086912284181518   0.3390208649613506   0.6245658180102851   0.9677781427256625   0.5339776078477825   0.1003217044772424
0.7242552944064735   0.25982216040053374   0.06927338914902487   0.5636510946754458   0.46616310699633245   0.4805265541207876   0.9699185064317586   0.5133272658641522   0.11053000791516347   0.42259643281100245   0.982613956687521   0.06233359376291303   0.054158516998731206   0.31591461591133   0.9425837041372624   0.21847928001111608   0.03866779060560675   0.6884734502656669   0.5338924757191107   0.8794584150497655   0.4141019725953217   0.7206953075400043   0.9999148678713282   0.7791367105725231   0.6898466781888482   0.46087314713947053   0.9306414787223033   0.2154856158970773   0.22368357119251572   0.980346593018683   0.9607229722905448   0.702158350032925   0.11315356327735225   0.5577501602076805   0.9781090156030238   0.639824756270012   0.058995046278621045   0.24183554429635049   0.03552531146576126   0.42134547625889596   0.02032725567301429   0.5533620940306836   0.5016328357466506   0.5418870612091304   0.6062252830776926   0.8326667864906794   0.5017179678753224   0.7627503506366075   0.9163786048888444   0.3717936393512088   0.5710764891530191   0.5472647347395301   0.6926950336963287   0.39144704633252586   0.6103535168624743   0.845106384706605   0.5795414704189764   0.8336968861248454   0.6322445012594506   0.20528162843659303   0.5205464241403553   0.5918613418284949   0.5967191897936893   0.7839361521776971
0.500219168467341   0.03849924779781124   0.09508635404703873   0.2420490909685666   0.8939938853896485   0.20583246130713193   0.5933683861717163   0.4792987403319592   0.9776152805008042   0.8340388219559232   0.022291897018697177   0.9320340055924291   0.2849202468044754   0.4425917756233973   0.41193838015622286   0.08692762088582404   0.7053787763854991   0.608894889498552   0.7796938788967722   0.881645992449231   0.18483235224514366   0.017033547670057072   0.1829746891030829   0.09770984027153393   0.6846131837778026   0.9785342998722458   0.08788833505604417   0.8556607493029673   0.790619298388154   0.7727018385651139   0.4945199488843279   0.37636200897100813   0.81300401788735   0.9386630166091908   0.4722280518656307   0.44432800337857903   0.5280837710828745   0.49607124098579347   0.060289671709407855   0.357400382492755   0.8227049946973756   0.8871763514872415   0.28059579281263564   0.475754390043524   0.6378726424522319   0.8701428038171845   0.09762110370955274   0.3780445497719901   0.9532594586744293   0.8916085039449386   0.009732768653508571   0.5223838004690228   0.16264016028627523   0.11890666537982474   0.5152128197691807   0.1460217914980146   0.34963614239892526   0.18024364877063395   0.042984767903550006   0.7016937881194356   0.8215523713160507   0.6841724077848405   0.9826950961941422   0.34429340562668054
0.9988473766186752   0.796996056297599   0.7020993033815065   0.8685390155831565   0.3609747341664433   0.9268532524804144   0.6044781996719538   0.49049446581116646   0.40771527549201403   0.03524474853547579   0.5947454310184452   0.9681106653421437   0.24507511520573882   0.916338083155651   0.07953261124926451   0.8220888738441291   0.8954389728068135   0.7360944343850171   0.03654784334571451   0.12039508572469354   0.07388660149076283   0.051922026600176634   0.05385274715157236   0.7761016800980131   0.07503922487208761   0.25492597030257774   0.35175344377006584   0.9075626645148565   0.7140644907056443   0.3280727178221633   0.7472752440981121   0.41706819870369   0.30634921521363023   0.2928279692866875   0.15252981307966682   0.4489575333615463   0.061274100007891415   0.37648988613103646   0.0729972018304023   0.6268686595174172   0.16583512720107785   0.6403954517460193   0.0364493584846878   0.5064735737927236   0.09194852571031503   0.5884734251458427   0.9825966113331155   0.7303718936947107   0.01690930083822742   0.333547454843265   0.6308431675630496   0.8228092291798542   0.30284481013258313   0.005474737021101704   0.8835679234649375   0.40574103047616417   0.9964955949189529   0.7126467677344142   0.7310381103852708   0.9567834971146179   0.9352214949110615   0.33615688160337776   0.6580409085548684   0.32991483759720064
0.7693863677099837   0.6957614298573584   0.6215915500701806   0.823441263804477   0.6774378419996686   0.10728800471151569   0.6389949387370651   0.09306937010976636   0.6605285411614412   0.7737405498682507   0.008151771174015596   0.2702601409299122   0.35768373102885803   0.768265812847149   0.12458384770907804   0.8645191104537481   0.36118813610990513   0.05561904511273479   0.3935457373238073   0.9077356133391302   0.4259666411988436   0.719462163509357   0.7355048287689389   0.5778207757419295   0.65658027348886   0.02370073365199863   0.11391327869875825   0.7543795119374526   0.9791424314891913   0.916412728940483   0.4749183399616931   0.6613101418276861   0.3186138903277501   0.14267217907223223   0.46676656878767747   0.391050000897774   0.960930159298892   0.3744063662250832   0.34218272107859943   0.5265308904440259   0.599742023188987   0.3187873211123485   0.9486369837547921   0.6187952771048958   0.17377538199014333   0.5993251576029914   0.21313215498585322   0.04097450136296624   0.5171951085012834   0.5756244239509928   0.09921887628709497   0.2865949894255137   0.538052677012092   0.6592116950105098   0.624300536325402   0.6252848475978275   0.21943878668434194   0.5165395159382776   0.15753396753772445   0.2342348467000536   0.2585086273854499   0.14213314971319435   0.815351246459125   0.7077039562560277
0.6587666041964629   0.8233458286008459   0.8667142627043329   0.0889086791511319   0.48499122220631957   0.2240206709978545   0.6535821077184797   0.047934177788165666   0.9677961137050362   0.6483962470468617   0.5543632314313847   0.7613391883626519   0.42974343669294407   0.9891845520363519   0.9300626951059828   0.13605434076482437   0.21030465000860216   0.4726450360980743   0.7725287275682583   0.9018194940647708   0.9517960226231523   0.33051188638487994   0.9571774811091334   0.1941155378087431   0.2930294184266894   0.507166057784034   0.0904632184048004   0.1052068586576112   0.8080381962203698   0.2831453867861795   0.43688111068632074   0.057272680869445536   0.8402420825153336   0.6347491397393178   0.8825178792549361   0.29593349250679357   0.41049864582238954   0.6455645877029659   0.9524551841489532   0.1598791517419692   0.2001939958137874   0.17291955160489164   0.17992645658069492   0.25805965767719846   0.2483979731906351   0.8424076652200118   0.2227489754715616   0.06394411986845534   0.9553685547639458   0.3352416074359777   0.1322857570667612   0.9587372612108441   0.14733035854357593   0.052096220649798214   0.6954046463804404   0.9014645803413986   0.3070882760282423   0.41734708091048045   0.8128867671255045   0.605531087834605   0.8965896302058527   0.7717824932075146   0.8604315829765512   0.4456519360926358
0.6963956343920653   0.5988629416026229   0.6805051263958563   0.18759227841543735   0.4479976612014302   0.7564552763826111   0.45775615092429467   0.12364815854698201   0.4926291064374845   0.4212136689466334   0.32547039385753346   0.16491089733613787   0.3452987478939086   0.36911744829683524   0.630065747477093   0.26344631699473925   0.038210471865666285   0.9517703673863548   0.8171789803515885   0.6579152291601342   0.14162084165981356   0.17998787417884027   0.9567473973750373   0.21226329306749847   0.4452252072677483   0.5811249325762173   0.2762422709791811   0.024671014652061115   0.997227546066318   0.8246696561936062   0.8184861200548864   0.9010228561050792   0.5045984396288336   0.4034559872469728   0.493015726197353   0.7361119587689412   0.15929969173492503   0.03433853895013757   0.86294997872026   0.472665641774202   0.12108921986925876   0.08256817156378277   0.045770998368671524   0.8147504126140678   0.9794683782094452   0.9025802973849425   0.08902360099363417   0.6024871195465693   0.5342431709416969   0.3214553648087251   0.8127813300144531   0.5778161048945082   0.5370156248753789   0.4967857086151189   0.9942952099595667   0.676793248789429   0.03241718524654527   0.0933297213681461   0.5012794837622137   0.9406812900204878   0.8731174935116203   0.058991182418008534   0.6383295050419535   0.46801564824628583
0.7520282736423615   0.9764230108542258   0.592558506673282   0.653265235632218   0.7725598954329163   0.07384271346928327   0.5035349056796479   0.05077811608564883   0.23831672449121938   0.7523873486605581   0.6907535756651948   0.4729620111911407   0.7013010996158405   0.2556016400454393   0.6964583657056281   0.7961687624017116   0.6688839143692953   0.16227191867729315   0.19517888194341457   0.8554874723812238   0.795766420857675   0.10328073625928462   0.5568493769014611   0.387471824134938   0.043738147215313515   0.12685772540505885   0.964290870228179   0.7342065885027199   0.27117825178239724   0.0530150119357756   0.4607559645485311   0.683428472417071   0.03286152729117785   0.30062766327521745   0.7700023888833364   0.21046646122593043   0.33156042767533733   0.04502602322977819   0.0735440231777082   0.4142976988242188   0.6626765133060422   0.882754104552485   0.8783651412342937   0.5588102264429949   0.8669100924483671   0.7794733682932004   0.3215157643328326   0.17133840230805691   0.8231719452330536   0.6526156428881416   0.3572248941046536   0.43713181380533694   0.5519936934506564   0.5996006309523659   0.8964689295561225   0.7537033413882659   0.5191321661594785   0.2989729676771485   0.1264665406727861   0.5432368801623354   0.1875717384841412   0.2539469444473703   0.0529225174950779   0.12893918133811666
0.5248952251780991   0.3711928398948853   0.17455737626078427   0.5701289548951217   0.6579851327297319   0.5917194716016849   0.8530416119279517   0.3987905525870648   0.8348131874966784   0.9391038287135434   0.49581671782329806   0.9616587387817278   0.282819494046022   0.3395031977611774   0.5993477882671756   0.207955397393462   0.7636873278865435   0.04053023008402891   0.47288124759438954   0.6647185172311265   0.5761155894024023   0.7865832856366586   0.4199587300993116   0.5357793358930099   0.05122036422430324   0.4153904457417733   0.24540135383852738   0.9656503809978881   0.3932352314945713   0.8236709741400885   0.3923597419105757   0.5668598284108234   0.5584220439978929   0.8845671454265451   0.8965430240872776   0.6052010896290955   0.2756025499518709   0.5450639476653677   0.297195235820102   0.3972456922356335   0.5119152220653274   0.5045337175813388   0.8243139882257124   0.7325271750045069   0.9357996326629251   0.7179504319446802   0.40435525812640083   0.19674783911149704   0.8845792684386218   0.30255998620290686   0.15895390428787348   0.23109745811360888   0.49134403694405054   0.4788890120628184   0.7665941623772978   0.6642376297027855   0.9329219929461576   0.5943218666362733   0.8700511382900201   0.059036540073690066   0.6573194429942868   0.049257918970905576   0.5728559024699181   0.6617908478380565
0.1454042209289594   0.5447242013895668   0.7485419142442057   0.9292636728335496   0.20960458826603434   0.8267737694448866   0.34418665611780486   0.7325158337220525   0.3250253198274125   0.5242137832419796   0.18523275182993135   0.5014183756084437   0.833681282883362   0.045324771179161234   0.41863858945263355   0.8371807459056582   0.9007592899372042   0.45100290454288794   0.5485874511626134   0.7781442058319681   0.24343984694291748   0.40174498557198235   0.9757315486926952   0.1163533579939115   0.09803562601395807   0.8570207841824156   0.22718963444848952   0.18708968516036187   0.8884310377479238   0.030247014737529068   0.8830029783306848   0.4545738514383093   0.5634057179205112   0.5060332314955495   0.6977702265007534   0.9531554758298656   0.7297244350371493   0.4607084603163882   0.27913163704811983   0.11597472992420746   0.828965145099945   0.009705555773500235   0.7305441858855064   0.3378305240922394   0.5855252981570276   0.6079605702015178   0.7548126371928112   0.22147716609832788   0.4874896721430695   0.7509397860191023   0.5276230027443217   0.03438748093796601   0.5990586343951457   0.7206927712815732   0.644620024413637   0.5798136294996568   0.035652916474634526   0.21465953978602378   0.9468497979128836   0.6266581536697912   0.30592848143748524   0.7539510794696356   0.6677181608647639   0.5106834237455836
0.4769633363375402   0.7442455236961354   0.9371739749792574   0.17285289965334427   0.8914380381805127   0.1362849534946175   0.18236133778644617   0.9513757335550164   0.40394836603744316   0.3853451674755152   0.6547383350421245   0.9169882526170504   0.8048897316422974   0.664652396193942   0.010118310628487497   0.33717462311739366   0.7692368151676628   0.44999285640791825   0.06326851271560387   0.7105164694476026   0.46330833373017766   0.6960417769382826   0.39555035185084003   0.1998330457020189   0.9863449973926375   0.9517962532421473   0.4583763768715826   0.026980146048674644   0.09490695921212479   0.8155112997475298   0.27601503908513647   0.07560441249365825   0.6909585931746817   0.43016613227201456   0.6212767040430119   0.15861615987660788   0.8860688615323842   0.7655137360780725   0.6111583934145245   0.8214415367592142   0.11683204636472135   0.31552087967015424   0.5478898806989206   0.11092506731161164   0.6535237126345437   0.6194791027318716   0.15233952884808058   0.9110920216095927   0.6671787152419063   0.6676828494897243   0.6939631519764979   0.8841118755609181   0.5722717560297815   0.8521715497421944   0.41794811289136147   0.8085074630672598   0.8813131628550999   0.42200541747017994   0.7966714088483495   0.6498913031906519   0.9952443013227156   0.6564916813921075   0.18551301543382503   0.8284497664314378
0.8784122549579942   0.3409708017219532   0.6376231347349044   0.7175246991198261   0.22488854232345057   0.7214916989900816   0.48528360588682384   0.8064326775102334   0.5577098270815443   0.05380884950035734   0.7913204539103259   0.9223208019493153   0.9854380710517628   0.20163729975816283   0.37337234101896444   0.11381333888205547   0.10412490819666298   0.7796318822879829   0.5767009321706149   0.4639220356914035   0.10888060687394735   0.12314020089587545   0.3911879167367899   0.6354722692599657   0.23046835191595308   0.7821693991739223   0.7535647820018855   0.9179475701401396   0.0055798095925025   0.06067770018384061   0.2682811761150616   0.11151489262990624   0.4478699825109582   0.006868850683483272   0.4769607222047357   0.18919409068059095   0.4624319114591954   0.8052315509253204   0.10358838118577128   0.07538075179853548   0.3583070032625324   0.02559966863733754   0.5268874490151564   0.611458716107132   0.24942639638858505   0.9024594677414621   0.13569953227836654   0.9759864468471662   0.01895804447263197   0.12029006856753985   0.3821347502764811   0.05803887670702659   0.01337823488012947   0.05961236838369924   0.11385357416141949   0.9465239840771204   0.5655082523691712   0.052743517700215965   0.6368928519566838   0.7573298933965295   0.1030763409099759   0.24751196677489554   0.5333044707709125   0.6819491415979939
0.7447693376474435   0.221912298137558   0.006417021755756116   0.07049042549086194   0.49534294125885847   0.3194528303960959   0.8707174894773896   0.09450397864369572   0.47638489678622653   0.19916276182855605   0.4885827392009085   0.03646510193666913   0.463006661906097   0.1395503934448568   0.374729165039489   0.08994111785954878   0.8974984095369257   0.08680687574464084   0.7378363130828052   0.3326112244630194   0.7944220686269499   0.8392949089697453   0.20453184231189273   0.6506620828650255   0.049652730979506336   0.6173826108321873   0.1981148205561366   0.5801716573741635   0.5543097897206478   0.2979297804360914   0.327397331078747   0.4856676787304678   0.07792489293442136   0.09876701860753535   0.8388145918778385   0.44920257679379866   0.6149182310283243   0.9592166251626786   0.4640854268383495   0.3592614589342499   0.7174198214913986   0.8724097494180377   0.7262491137555442   0.026650234471230508   0.9229977528644487   0.03311484044829239   0.5217172714436515   0.375988151606205   0.8733450218849423   0.41573222961610506   0.32360245088751494   0.7958164942320415   0.3190352321642945   0.11780244918001367   0.9962051198087679   0.3101488155015737   0.24111033922987316   0.019035430572478324   0.15739052793092942   0.8609462387077751   0.6261921082015488   0.05981880540979978   0.6933051010925799   0.5016847797735252
0.9087722867101503   0.18740905599176208   0.9670559873370357   0.47503454530229466   0.9857745338457016   0.1542942155434697   0.4453387158933841   0.09904639369608961   0.11242951196075919   0.7385619859273647   0.12173626500586915   0.3032298994640481   0.7933942797964647   0.620759536747351   0.12553114519710123   0.9930810839624744   0.5522839405665915   0.6017241061748726   0.9681406172661718   0.13213484525469932   0.9260918323650427   0.5419053007650728   0.27483551617359187   0.6304500654811741   0.01731954565489237   0.35449624477331076   0.30777952883655624   0.1554155201788795   0.0315450118091908   0.20020202922984107   0.8624408129431721   0.0563691264827899   0.9191154998484317   0.46164004330247643   0.740704547937303   0.7531392270187418   0.12572122005196695   0.8408805065551255   0.6151734027402017   0.7600581430562674   0.5734372794853755   0.23915640038025288   0.64703278547403   0.6279232978015681   0.6473454471203328   0.6972510996151801   0.37219726930043806   0.997473232320394   0.6300259014654405   0.3427548548418693   0.06441774046388182   0.8420577121415145   0.5984808896562496   0.14255282561202823   0.2019769275207097   0.7856885856587246   0.679365389807818   0.6809127823095518   0.4612723795834067   0.032549358639982755   0.5536441697558511   0.8400322757544263   0.8460989768432049   0.2724912155837153
0.9802068902704756   0.6008758753741734   0.199066191369175   0.6445679177821472   0.33286144315014277   0.9036247757589934   0.826868922068737   0.6470946854617532   0.7028355416847024   0.5608699209171241   0.7624511816048551   0.8050369733202387   0.10435465202845273   0.41831709530509587   0.5604742540841454   0.019348387661514196   0.4249892622206347   0.7374043129955441   0.0992018745007387   0.9867990290215315   0.8713450924647836   0.8973720372411178   0.25310289765753374   0.7143078134378161   0.8911382021943081   0.29649616186694433   0.054036706288358764   0.06973989565566895   0.5582767590441653   0.3928713861079509   0.22716778421962183   0.4226452101939157   0.855441217359463   0.8320014651908268   0.4647166026147667   0.6176082368736769   0.7510865653310101   0.413684369885731   0.9042423485306214   0.5982598492121628   0.3260973031103755   0.6762800568901869   0.8050404740298827   0.6114608201906313   0.4547522106455918   0.7789080196490692   0.5519375763723489   0.8971530067528152   0.5636140084512837   0.48241185778212486   0.4979008700839901   0.8274131110971462   0.005337249407118401   0.08954047167417391   0.2707330858643683   0.4047679009032305   0.14989603204765548   0.2575390064833471   0.8060164832496015   0.7871596640295535   0.39880946671664524   0.8438546365976161   0.9017741347189802   0.18889981481739077
0.0727121636062698   0.16757457970742917   0.09673366068909756   0.5774389946267594   0.617959952960678   0.38866656005836   0.5447960843167486   0.6802859878739442   0.05434594450939431   0.9062547022762352   0.04689521423275858   0.852872876776798   0.04900869510227591   0.8167142306020613   0.7761621283683903   0.44810497587356746   0.8991126630546205   0.5591752241187141   0.9701456451187888   0.660945311844014   0.5003031963379752   0.7153205875210981   0.0683715103998086   0.47204549702662313   0.4275910327317054   0.5477460078136689   0.971637849710711   0.8946065023998637   0.8096310797710273   0.15907944775530888   0.42684176539396235   0.2143205145259195   0.7552851352616331   0.25282474547907374   0.3799465511612038   0.36144763774912153   0.7062764401593572   0.4361105148770125   0.6037844227928134   0.913342661875554   0.8071637771047367   0.8769352907582983   0.6336387776740247   0.2523973500315401   0.30686058076676154   0.16161470323720026   0.5652672672742161   0.7803518530049169   0.8792695480350562   0.6138686954235314   0.5936294175635051   0.8857453506050533   0.06963846826402877   0.4547892476682225   0.1667876521695427   0.6714248360791338   0.3143533330023957   0.20196450218914874   0.7868411010083389   0.30997719833001225   0.6080768928430386   0.7658539873121363   0.18305667821552546   0.39663453645445823
0.8009131157383018   0.8889186965538379   0.5494179005415007   0.14423718642291808   0.49405253497154034   0.7273039933166376   0.9841506332672847   0.3638853334180011   0.6147829869364841   0.11343529789310627   0.3905212157037797   0.47813998281294784   0.5451445186724554   0.6586460502248838   0.22373356353423698   0.8067151467338141   0.23079118567005968   0.456681548035735   0.4368924625258981   0.49673794840380175   0.6227142928270212   0.6908275607235989   0.2538357843103726   0.10010341194934354   0.8218011770887192   0.8019088641697609   0.7044178837688718   0.9558662255264254   0.32774864211717897   0.07460487085312326   0.7202672505015871   0.5919808921084243   0.7129656551806948   0.961169572960017   0.3297460347978074   0.11384090929547654   0.1678211365082394   0.3025235227351332   0.10601247126357043   0.3071257625616625   0.9370299508381797   0.8458419746993981   0.6691200087376724   0.8103878141578608   0.31431565801115857   0.15501441397579935   0.4152842244272998   0.7102844022085172   0.4925144809224393   0.3531055498060385   0.7108663406584279   0.7544181766820918   0.16476583880526033   0.2785006789529152   0.9905990901568409   0.16243728457366738   0.45180018362456553   0.3173311059928982   0.6608530553590335   0.04859637527819084   0.2839790471163261   0.014807583257765013   0.554840584095463   0.7414706127165284
0.34694909627814635   0.16896560855836687   0.8857205753577907   0.9310827985586676   0.03263343826698777   0.013951194582567503   0.4704363509304909   0.22079839635015042   0.5401189573445485   0.6608456447765291   0.759570010272063   0.4663802196680587   0.37535311853928816   0.3823449658236138   0.7689709201152221   0.3039429350943913   0.9235529349147227   0.06501385983071563   0.10811786475618865   0.25534655981620047   0.6395738877983965   0.05020627657295062   0.5532772806607256   0.5138759470996721   0.29262479152025017   0.8812406680145838   0.667556705302935   0.5827931485410045   0.2599913532532624   0.8672894734320162   0.19712035437244405   0.3619947521908541   0.719872395908714   0.20644382865548722   0.4375503441003811   0.8956145325227953   0.3445192773694258   0.8240988628318734   0.668579423985159   0.591671597428404   0.4209663424547031   0.7590850030011578   0.5604615592289703   0.3363250376122036   0.7813924546563066   0.7088787264282072   0.007184278568244732   0.8224490905125315   0.48876766313605635   0.8276380584136234   0.3396275732653098   0.23965594197152698   0.22877630988279396   0.9603485849816071   0.14250721889286574   0.8776611897806729   0.50890391397408   0.7539047563261199   0.7049568747924847   0.9820466572578775   0.16438463660465424   0.9298058934942466   0.03637745080732568   0.3903750598294735
0.7434182941499511   0.17072089049308878   0.47591589157835534   0.05405002221726989   0.9620258394936445   0.46184216406488166   0.4687316130101106   0.23160093170473842   0.47325817635758816   0.6342041056512583   0.1291040397448008   0.9919449897332114   0.2444818664747942   0.6738555206696512   0.9865968208519351   0.11428379995253851   0.7355779525007142   0.9199507643435313   0.2816399460594504   0.13223714269466097   0.5711933158960599   0.9901448708492848   0.2452624952521247   0.7418620828651875   0.8277750217461088   0.819423980356196   0.7693466036737694   0.6878120606479176   0.8657491822524643   0.3575818162913143   0.30061499066365877   0.45621112894317917   0.3924910058948762   0.7233777106400561   0.17151095091885796   0.46426613920996773   0.14800913942008195   0.04952218997040481   0.1849141300669229   0.3499823392574292   0.41243118691936775   0.12957142562687352   0.9032741840074725   0.21774519656276828   0.8412378710233078   0.13942655477758872   0.6580116887553478   0.4758831136975808   0.013462849277198954   0.32000257442139274   0.8886650850815784   0.7880710530496632   0.14771366702473462   0.9624207581300784   0.5880500944179197   0.33185992410648407   0.7552226611298585   0.2390430474900224   0.4165391434990616   0.8675937848965163   0.6072135217097765   0.18952085751961759   0.23162501343213873   0.5176114456390871
0.1947823347904087   0.05994943189274408   0.32835082942466626   0.2998662490763188   0.3535444637671009   0.9205228771151553   0.6703391406693184   0.823983135378738   0.34008161448990193   0.6005203026937627   0.7816740555877401   0.035912082329074765   0.19236794746516733   0.6380995445636842   0.19362396116982042   0.7040521582225907   0.43714528633530886   0.3990564970736618   0.7770848176707588   0.8364583733260744   0.8299317646255324   0.2095356395540442   0.5454598042386201   0.3188469276869873   0.6351494298351237   0.14958620766130012   0.2171089748139538   0.0189806786106685   0.28160496606802277   0.22906333054614478   0.5467698341446353   0.1949975432319305   0.9415233515781208   0.6285430278523821   0.7650957785568953   0.15908546090285575   0.7491554041129534   0.990443483288698   0.5714718173870749   0.45503330268026504   0.3120101177776446   0.5913869862150362   0.7943869997163161   0.6185749293541907   0.4820783531521122   0.38185134666099196   0.24892719547769607   0.29972800166720337   0.8469289233169885   0.23226513899969184   0.03181822066374228   0.2807473230565348   0.5653239572489658   0.0032018084535470745   0.4850483865191069   0.08574977982460434   0.623800605670845   0.3746587806011649   0.7199526079622116   0.9266643189217486   0.8746452015578915   0.38421529731246695   0.14848079057513675   0.47163101624148357
0.562635083780247   0.7928283110974308   0.35409379085882065   0.853056086887293   0.08055673062813468   0.4109769644364388   0.10516659538112455   0.5533280852200896   0.2336278073111461   0.1787118254367469   0.07334837471738227   0.2725807621635547   0.6683038500621803   0.17551001698319985   0.5882999881982753   0.18683098233895037   0.044503244391335295   0.8008512363820349   0.8683473802360637   0.2601666634172018   0.16985804283344377   0.41663593906956803   0.719866589660927   0.7885356471757182   0.6072229590531969   0.6238076279721373   0.36577279880210634   0.9354795602884253   0.5266662284250622   0.2128306635356985   0.2606062034209818   0.3821514750683357   0.2930384211139161   0.03411883809895157   0.18725782870359953   0.10957071290478097   0.6247345710517358   0.8586088211157518   0.5989578405053242   0.9227397305658306   0.5802313266604004   0.05775758473371679   0.7306104602692605   0.6625730671486288   0.4103732838269567   0.6411216456641488   0.010743870608333471   0.8740374199729106   0.8031503247737598   0.01731401769201153   0.6449710718062271   0.9385578596844854   0.2764840963486977   0.804483354156313   0.3843648683852453   0.5564063846161497   0.9834456752347815   0.7703645160573614   0.19710703968164578   0.4468356717113687   0.3587111041830458   0.9117556949416098   0.5981491991763216   0.5240959411455381
0.7784797775226453   0.853998110207893   0.8675387389070611   0.8615228739969093   0.3681064936956886   0.21287646454374418   0.8567948682987276   0.9874854540239987   0.5649561689219288   0.19556244685173266   0.21182379649250055   0.04892759433951329   0.2884720725732311   0.39107909269541963   0.8274589281072553   0.4925212097233636   0.3050263973384495   0.6207145766380582   0.6303518884256094   0.045685538011994924   0.9463152931554036   0.7089588816964484   0.032202689249287854   0.5215895968664568   0.16783551563275834   0.8549607714885554   0.1646639503422267   0.6600667228695475   0.7997290219370697   0.6420843069448112   0.30786908204349905   0.6725812688455489   0.23477285301514095   0.4465218600930786   0.09604528555099848   0.6236536745060356   0.9463007804419099   0.055442767397659014   0.2685863574437432   0.131132464782672   0.6412743831034604   0.4347281907596009   0.6382344690181337   0.08544692677067706   0.6949590899480568   0.7257693090631525   0.6060317797688459   0.5638573299042202   0.5271235743152984   0.8708085375745971   0.44136782942661923   0.9037906070346727   0.7273945523782287   0.2287242306297858   0.13349874738312018   0.23120933818912381   0.49262169936308775   0.7822023705367072   0.037453461832121705   0.6075556636830882   0.5463209189211778   0.7267596031390482   0.7688671043883785   0.47642319890041623
0.9050465358177174   0.2920314123794473   0.13063263537024472   0.3909762721297392   0.21008744586966074   0.5662621033162948   0.5246008556013988   0.827118942225519   0.6829638715543623   0.6954535657416977   0.0832330261747796   0.9233283351908462   0.9555693191761336   0.46672933511191195   0.9497342787916594   0.6921189970017224   0.4629476198130459   0.6845269645752048   0.9122808169595377   0.0845633333186342   0.916626700891868   0.9577673614361566   0.14341371257115923   0.6081401344182179   0.011580165074150515   0.6657359490567093   0.012781077200914528   0.21716386228847875   0.8014927192044897   0.09947384574041446   0.48818022159951574   0.3900449200629598   0.11852884765012744   0.4040202799987167   0.4049471954247361   0.46671658487211354   0.1629595284739938   0.9372909448868048   0.4552129166330767   0.7745975878703911   0.700011908660948   0.2527639803116   0.5429320996735391   0.6900342545517569   0.7833852077690799   0.2949966188754435   0.39951838710237975   0.08189412013353896   0.7718050426949294   0.6292606698187342   0.38673730990146526   0.8647302578450602   0.9703123234904396   0.5297868240783198   0.8985570883019495   0.4746853377821004   0.8517834758403122   0.12576654407960303   0.49360989287721335   0.007968752909986864   0.6888239473663184   0.18847559919279824   0.03839697624413665   0.23337116503959573
0.9888120387053705   0.9357116188811982   0.4954648765705976   0.5433369104878388   0.2054268309362905   0.6407150000057548   0.09594648946821786   0.46144279035429986   0.43362178824136105   0.011454330187020561   0.7092091795667527   0.5967125325092396   0.4633094647509214   0.48166750610870085   0.8106520912648031   0.12202719472713924   0.6115259889106092   0.3559009620290978   0.31704219838758974   0.11405844181715238   0.9227020415442908   0.16742536283629958   0.2786452221434531   0.8806872767775566   0.9338900028389203   0.23171374395510136   0.7831803455728554   0.3373503662897178   0.7284631719026299   0.5909987439493466   0.6872338561046376   0.8759075759354179   0.2948413836612688   0.579544413762326   0.9780246765378849   0.2791950434261783   0.8315319189103474   0.09787690765362521   0.16737258527308185   0.15716784869903902   0.22000592999973817   0.7419759456245274   0.8503303868854921   0.043109406881886636   0.29730388845544736   0.5745505827882278   0.571685164742039   0.16242213010433001   0.36341388561652704   0.3428368388331265   0.7885048191691835   0.8250717638146122   0.6349507137138972   0.7518380948837798   0.10127096306454592   0.9491641878791942   0.34010933005262844   0.17229368112145385   0.12324628652666095   0.669969144453016   0.508577411142281   0.07441677346782864   0.9558737012535791   0.5128012957539769
0.28857148114254294   0.33244082784330126   0.105543314368087   0.46969188887209035   0.9912675926870955   0.7578902450550734   0.533858149626048   0.3072697587677603   0.6278537070705685   0.4150534062219469   0.7453533304568645   0.48219799495314813   0.9929029933566713   0.663215311338167   0.6440823673923186   0.5330338070739539   0.6527936633040429   0.4909216302167132   0.5208360808656576   0.8630646626209378   0.1442162521617618   0.41650485674888454   0.5649623796120785   0.3502633668669609   0.8556447710192189   0.08406402890558332   0.4594190652439915   0.8805714779948706   0.8643771783321232   0.32617378385050994   0.9255609156179435   0.5733017192271103   0.23652347126155474   0.911120377628563   0.18020758516107901   0.09110372427396216   0.2436204779048834   0.24790506629039596   0.5361252177687604   0.5580699172000083   0.5908268146008405   0.7569834360736828   0.01528913690310281   0.6950052545790704   0.4466105624390787   0.34047857932479825   0.4503267572910243   0.3447418877121095   0.5909657914198598   0.2564145504192149   0.9909076920470328   0.4641704097172389   0.7265886130877366   0.930240766568705   0.06534677642908925   0.8908686904901286   0.4900651418261818   0.01912038894014201   0.8851391912680102   0.7997649662161664   0.24644466392129843   0.771215322649746   0.3490139734992498   0.24169504901615818
0.655617849320458   0.014231886576063271   0.333724836596147   0.5466897944370878   0.20900728688137923   0.673753307251265   0.8833980793051227   0.20194790672497828   0.6180414954615194   0.41733875683205013   0.8924903872580899   0.7377774970077394   0.8914528823737828   0.4870979902633451   0.8271436108290007   0.8469088065176108   0.401387740547601   0.4679776013232031   0.9420044195609905   0.04714384030144429   0.15494307662630258   0.6967622786734571   0.5929904460617407   0.8054487912852861   0.49932522730584467   0.6825303920973937   0.25926560946559374   0.25875899684819836   0.2903179404244654   0.008777084846128744   0.37586753016047103   0.05681109012322008   0.672276444962946   0.5914383280140786   0.4833771429023811   0.3190335931154807   0.7808235625891632   0.10434033775073351   0.6562335320733804   0.47212478659786994   0.3794358220415621   0.6363627364275304   0.7142291125123899   0.42498094629642563   0.22449274541525957   0.9396004577540733   0.12123866645064921   0.6195321550111396   0.7251675181094149   0.25707006565667956   0.8619730569850554   0.3607731581629412   0.43484957768494953   0.24829298081055082   0.48610552682458447   0.3039620680397211   0.7625731327220036   0.6568546527964721   0.002728383922203403   0.9849284749242404   0.9817495701328404   0.5525143150457387   0.346494851848823   0.5128036883263705
0.6023137480912782   0.9161515786182083   0.6322657393364332   0.08782274202994478   0.37782100267601865   0.976551120864135   0.511027072885784   0.46829058701880527   0.6526534845666037   0.7194810552074554   0.6490540159007284   0.10751742885586407   0.21780390688165419   0.4711880743969046   0.16294848907614395   0.803555360816143   0.4552307741596507   0.8143334216004324   0.16022010515394053   0.8186268858919026   0.4734812040268103   0.2618191065546937   0.8137252533051175   0.30582319756553217   0.8711674559355321   0.3456675279364854   0.18145951396868437   0.21800045553558736   0.49334645325951354   0.36911640707235044   0.6704324410829005   0.7497098685167821   0.8406929686929098   0.6496353518648951   0.02137842518217204   0.642192439660918   0.6228890618112556   0.17844727746799052   0.8584299361060281   0.8386370788447751   0.16765828765160493   0.3641138558675581   0.6982098309520876   0.020010192952872482   0.6941770836247946   0.10229474931286446   0.8844845776469701   0.7141869953873403   0.8230096276892624   0.756627221376379   0.7030250636782857   0.496186539851753   0.3296631744297489   0.38751081430402856   0.0325926225953852   0.7464766713349709   0.4889702057368391   0.7378754624391335   0.011214197413213159   0.10428423167405282   0.8660811439255836   0.559428184971143   0.15278426130718506   0.26564715282927776
0.6984228562739786   0.19531432910358484   0.4545744303550975   0.24563695987640527   0.004245772649184017   0.09301957979072038   0.5700898527081274   0.5314499644890649   0.1812361449599216   0.33639235841434134   0.8670647890298417   0.03526342463731197   0.8515729705301727   0.9488815441103128   0.8344721664344565   0.2887867533023411   0.3626027647933336   0.21100608167117924   0.8232579690212434   0.18450252162828829   0.4965216208677501   0.6515778967000363   0.6704737077140583   0.9188553687990105   0.7980987645937715   0.4562635675964514   0.21589927735896086   0.6732184089226052   0.7938529919445875   0.36324398780573103   0.6458094246508335   0.1417684444335403   0.6126168469846659   0.026851629391389686   0.7787446356209916   0.10650501979622834   0.7610438764544932   0.07797008528107693   0.9442724691865351   0.8177182664938872   0.3984411116611596   0.8669640036098977   0.12101450016529161   0.633215744865599   0.9019194907934095   0.21538610690986143   0.45054079245123324   0.7143603760665884   0.10382072619963802   0.75912253931341   0.23464151509227238   0.041141967143983195   0.30996773425505053   0.395878551507679   0.5888320904414389   0.8993735227104429   0.6973508872703846   0.3690269221162893   0.8100874548204473   0.7928685029142145   0.9363070108158914   0.2910568368352124   0.8658149856339122   0.9751502364203273
0.5378658991547318   0.42409283322531466   0.7448004854686207   0.3419344915547284   0.6359464083613223   0.20870672631545326   0.2942596930173874   0.6275741154881399   0.5321256821616843   0.4495841870020432   0.05961817792511505   0.5864321483441567   0.2221579479066338   0.05370563549436423   0.47078608748367606   0.6870586256337138   0.5248070606362492   0.684678713378075   0.6606986326632287   0.8941901227194993   0.5885000498203578   0.39362187654286257   0.7948836470293165   0.919039886299172   0.050634150665625884   0.9695290433175479   0.050083161560695776   0.5771053947444436   0.41468774230430355   0.7608223170020947   0.7558234685433084   0.9495312792563037   0.8825620601426193   0.3112381300000514   0.6962052906181933   0.3630991309121469   0.6604041122359855   0.25753249450568716   0.22541920313451722   0.6760405052784331   0.13559705159973634   0.5728537811276122   0.5647205704712884   0.7818503825589338   0.5470970017793786   0.1792319045847497   0.7698369234419721   0.8628104962597618   0.49646285111375277   0.2097028612672018   0.7197537618812763   0.28570510151531825   0.08177510880944917   0.44888054426510715   0.9639302933379679   0.3361738222590146   0.1992130486668299   0.13764241426505577   0.2677250027197746   0.9730746913468676   0.5388089364308444   0.8801099197593686   0.042305799585257375   0.29703418606843457
0.4032118848311081   0.3072561386317563   0.4775852291139689   0.5151838035095008   0.8561148830517294   0.12802423404700664   0.7077483056719969   0.652373307249739   0.35965203193797673   0.9183213727798049   0.9879945437907206   0.36666820573442066   0.2778769231285275   0.46944082851469765   0.02406425045275273   0.03049438347540603   0.07866387446169763   0.33179841424964185   0.7563392477329781   0.05741969212853835   0.5398549380308532   0.4516884944902733   0.7140334481477207   0.7603855060601038   0.13664305319974512   0.14443235585851696   0.23644821903375185   0.245201702550603   0.2805281701480157   0.01640812181151034   0.528699913361755   0.5928283953008641   0.920876138210039   0.09808674903170553   0.5407053695710343   0.22616018956644343   0.6429992150815114   0.6286459205170079   0.5166411191182816   0.1956658060910374   0.5643353406198138   0.296847506267366   0.7603018713853035   0.13824611396249906   0.024480402588960577   0.8451590117770927   0.04626842323758274   0.3778606079023953   0.8878373493892154   0.7007266559185757   0.8098202042038308   0.1326589053517923   0.6073091792411998   0.6843185341070654   0.2811202908420759   0.5398305100509282   0.6864330410311608   0.5862317850753599   0.7404149212710416   0.3136703204844848   0.043433825949649396   0.957585864558352   0.2237738021527599   0.11800451439344739
0.4790984853298356   0.660738358290986   0.4634719307674564   0.9797584004309483   0.454618082740875   0.8155793465138933   0.4172035075298737   0.601897792528553   0.5667807333516596   0.1148526905953175   0.6073833033260427   0.4692388871767607   0.9594715541104598   0.43053415648825205   0.3262630124839669   0.9294083771258325   0.273038513079299   0.8443023714128922   0.5858480912129254   0.6157380566413477   0.2296046871296496   0.8867165068545402   0.3620742890601655   0.4977335422479003   0.750506201799814   0.22597814856355417   0.8986023582927091   0.5179751418169519   0.29588811905893897   0.41039880204966095   0.4813988507628354   0.9160773492883989   0.7291073857072794   0.29554611145434345   0.8740155474367927   0.4468384621116382   0.7696358315968196   0.8650119549660914   0.5477525349528257   0.5174300849858057   0.49659731851752054   0.020709583553199195   0.9619044437399004   0.901692028344458   0.26699263138787094   0.13399307669865904   0.5998301546797349   0.4039584860965577   0.516486429588057   0.9080149281351049   0.7012277963870258   0.8859833442796057   0.22059831052911802   0.4976161260854439   0.21982894562419045   0.9699059949912068   0.49149092482183865   0.2020700146311005   0.3458133981873978   0.5230675328795686   0.7218550932250191   0.3370580596650091   0.7980608632345721   0.0056374478937629025
0.22525777470749853   0.31634847611180994   0.8361564194946718   0.10394541954930489   0.9582651433196275   0.1823553994131509   0.23632626481493682   0.6999869334527472   0.4417787137315706   0.27434047127804606   0.535098468427911   0.8140035891731414   0.22118040320245258   0.7767243451926021   0.31526952280372056   0.8440975941819346   0.7296894783806139   0.5746543305615016   0.9694561246163227   0.32103006130236605   0.00783438515559487   0.2375962708964925   0.1713952613817506   0.31539261340860314   0.7825766104480963   0.9212477947846825   0.33523884188707886   0.21144719385929825   0.8243114671284688   0.7388923953715316   0.09891257707214203   0.511460260406551   0.3825327533968982   0.46455192409348556   0.5638141086442311   0.6974566712334096   0.16135235019444558   0.6878275789008834   0.2485445858405105   0.853359077051475   0.4316628718138316   0.11317324833938185   0.2790884612241878   0.5323290157491088   0.42382848665823675   0.8755769774428893   0.1076931998424372   0.21693640234050574   0.6412518762101405   0.9543291826582069   0.7724543579553583   0.0054892084812074825   0.8169404090816716   0.2154367872866752   0.6735417808832164   0.4940289480746564   0.43440765568477346   0.7508848631931896   0.10972767223898526   0.7965722768412469   0.27305530549032786   0.06305728429230614   0.8611830863984747   0.9432131997897719
0.8413924336764963   0.9498840359529243   0.5820946251742869   0.410884184040663   0.4175639470182595   0.07430705851003494   0.47440142533184976   0.19394778170015728   0.776312070808119   0.11997787585182812   0.7019470673764914   0.1884585732189498   0.9593716617264475   0.9045410885651529   0.028405286493275082   0.6944296251442934   0.524964006041674   0.15365622537196333   0.9186776142542898   0.8978573483030465   0.2519087005513461   0.09059894107965717   0.05749452785581506   0.9546441485132746   0.4105162668748498   0.14071490512673288   0.4753999026815281   0.5437599644726117   0.9929523198565904   0.06640784661669792   0.0009984773496783707   0.34981218277245435   0.21664024904847126   0.9464299707648698   0.29905140997318697   0.16135360955350456   0.2572685873220238   0.04188888219971687   0.2706461234799119   0.4669239844092112   0.7323045812803498   0.8882326568277535   0.35196850922562206   0.5690666361061647   0.48039588072900374   0.7976337157480964   0.294473981369807   0.61442248759289   0.0698796138541539   0.6569188106213635   0.8190740786882789   0.07066252312027839   0.07692729399756355   0.5905109640046656   0.8180756013386006   0.720850340347824   0.8602870449490922   0.6440809932397957   0.5190241913654136   0.5594967307943195   0.6030184576270685   0.602192111040079   0.24837806788550165   0.09257274638510826
0.8707138763467187   0.7139594542123253   0.8964095586598796   0.5235061102789436   0.39031799561771496   0.916325738464229   0.6019355772900726   0.9090836226860536   0.32043838176356104   0.2594069278428655   0.7828614986017937   0.8384210995657752   0.2435110877659975   0.6688959638381999   0.9647858972631932   0.11757075921795117   0.3832240428169052   0.02481497059840413   0.4457617058977796   0.5580740284236317   0.7802055851898367   0.42262285955832524   0.19738363801227793   0.4655012820385234   0.909491708843118   0.7086634053459998   0.30097407935239834   0.9419951717595798   0.5191737132254031   0.7923376668817709   0.6990385020623258   0.03291154907352625   0.19873533146184205   0.5329307390389053   0.9161770034605321   0.19449044950775105   0.9552242436958446   0.8640347752007055   0.9513911061973389   0.07691969028979988   0.5720002008789393   0.8392198046023013   0.5056294002995594   0.5188456618661682   0.7917946156891027   0.4165969450439761   0.3082457622872814   0.05334437982764473   0.8823029068459846   0.7079335396979762   0.007271682934883077   0.11134920806806489   0.3631291936205815   0.9155958728162054   0.3082331808725573   0.07843765899453864   0.1643938621587394   0.38266513377730005   0.39205617741202525   0.8839472094867876   0.20916961846289486   0.5186303585765946   0.4406650712146863   0.8070275191969877
0.6371694175839555   0.6794105539742933   0.935035670915127   0.2881818573308195   0.8453748018948528   0.2628136089303172   0.6267899086278456   0.2348374775031748   0.9630718950488683   0.554880069232341   0.6195182256929624   0.1234882694351099   0.5999427014282868   0.6392841964161355   0.31128504482040514   0.04505061044057128   0.43554883926954735   0.2566190626388355   0.91922886740838   0.1611034009537837   0.2263792208066525   0.7379887040622409   0.4785637961936936   0.354075881756796   0.589209803222697   0.05857815008794759   0.5435281252785666   0.06589402442597647   0.7438350013278442   0.7957645411576304   0.9167382166507211   0.8310565469228017   0.7807631062789759   0.24088447192528942   0.2972199909577586   0.7075682774876918   0.18082040485068915   0.6016002755091538   0.9859349461373534   0.6625176670471205   0.7452715655811418   0.34498121287031835   0.06670607872897351   0.5014142660933368   0.5188923447744893   0.6069925088080774   0.5881422825352799   0.14733838433654078   0.9296825415517923   0.5484143587201299   0.04461415725671326   0.08144435991056431   0.18584754022394817   0.7526498175624995   0.1278759406059922   0.25038781298776264   0.4050844339449723   0.5117653456372101   0.8306559496482336   0.5428195355000709   0.22426402909428314   0.9101650701280563   0.8447210035108802   0.8803018684529503
0.47899246351314134   0.5651838572577379   0.7780149247819066   0.3788876023596136   0.960100118738652   0.9581913484496604   0.18987264224662675   0.2315492180230728   0.03041757718685971   0.4097769897295305   0.14525848498991348   0.15010485811250848   0.8445700369629116   0.657127172167031   0.017382544383921304   0.8997170451247458   0.43948560301793926   0.14536182652982096   0.18672659473568773   0.356897509624675   0.21522157392365615   0.23519675640176477   0.34200559122480756   0.4765956411717246   0.7362291104105148   0.670012899144027   0.5639906664429009   0.09770803881211101   0.7761289916718628   0.7118215506943665   0.37411802419627416   0.8661588207890382   0.7457114144850031   0.302044560964836   0.22885953920636068   0.7160539626765298   0.9011413775220916   0.644917388797805   0.21147699482243937   0.8163369175517838   0.46165577450415224   0.49955556226798403   0.024750400086751657   0.4594394079271089   0.24643420058049612   0.2643588058662193   0.6827448088619441   0.9828437667553843   0.5102050901699813   0.5943459067221923   0.11875414241904318   0.8851357279432732   0.7340760984981185   0.8825243560278259   0.744636118222769   0.018976907154235067   0.9883646840131155   0.5804797950629899   0.5157765790164084   0.30292294447770535   0.08722330649102393   0.9355624062651848   0.30429958419396896   0.48658602692592146
0.6255675319868716   0.4360068439972008   0.2795491841072173   0.027146618998812596   0.37913333140637556   0.17164803813098153   0.5968043752452732   0.044302852243428316   0.8689282412363942   0.5773021314087892   0.47805023282623005   0.15916712430015503   0.13485214273827575   0.6947777753809633   0.733414114603461   0.14019021714591998   0.14648745872516028   0.11429798031797349   0.21763753558705265   0.8372672726682147   0.059264152234136364   0.17873557405278864   0.9133379513930837   0.35068124574229315   0.4336966202472647   0.7427287300555878   0.6337887672858664   0.32353462674348055   0.054563288840889124   0.5710806919246063   0.036984392040593145   0.2792317745000522   0.18563504760449487   0.9937785605158171   0.5589341592143631   0.12006465019989719   0.05078290486621912   0.29900078513485384   0.8255200446109021   0.9798744330539773   0.9042954461410588   0.18470280481688034   0.6078825090238494   0.1426071603857626   0.8450312939069224   0.005967230764091709   0.6945445576307657   0.7919259146434695   0.41133467365965776   0.26323850070850385   0.060755790344899405   0.4683912878999889   0.35677138481876863   0.6921578087838975   0.02377139830430626   0.18915951339993667   0.1711363372142738   0.6983792482680804   0.4648372390899431   0.06909486320003949   0.12035343234805466   0.3993784631332266   0.639317194479041   0.08922043014606226
0.21605798620699584   0.21467565831634625   0.031434685455191576   0.9466132697602997   0.37102669230007335   0.20870842755225452   0.3368901278244258   0.1546873551168302   0.9596920186404156   0.9454699268437506   0.27613433747952637   0.6862960672168413   0.602920633821647   0.2533121180598531   0.2523629391752201   0.49713655381690464   0.43178429660737316   0.5549328697917727   0.787525700085277   0.42804169061686514   0.31143086425931854   0.15555440665854608   0.14820850560623597   0.33882126047080285   0.09537287805232268   0.9408787483421999   0.11677382015104439   0.3922079907105032   0.7243461857522493   0.7321703207899454   0.7798836923266186   0.23752063559367298   0.7646541671118338   0.7867003939461946   0.5037493548470922   0.5512245683768316   0.16173353329018675   0.5333882758863416   0.25138641567187203   0.054088014559927074   0.7299492366828135   0.9784554060945689   0.4638607155865951   0.6260463239430619   0.41851837242349504   0.8229009994360228   0.3156522099803591   0.28722506347225907   0.32314549437117235   0.882022251093823   0.19887838982931472   0.8950170727617559   0.598799308618923   0.14985193030387767   0.41899469750269613   0.6574964371680829   0.8341451415070893   0.363151536357683   0.915245342655604   0.1062718687912512   0.6724116082169026   0.8297632604713414   0.663858926983732   0.052183854231324114
0.942462371534089   0.8513078543767725   0.19999821139713683   0.4261375302882622   0.523943999110594   0.028406854940749682   0.8843460014167778   0.1389124668160031   0.2007985047394216   0.1463846038469267   0.685467611587463   0.24389539405424723   0.6019991961204986   0.996532673543049   0.26647291408476687   0.5863989568861644   0.7678540546134093   0.633381137185366   0.35122757142916294   0.48012708809491317   0.09544244639650663   0.8036178767140246   0.687368644445431   0.427943233863589   0.15298007486241763   0.952310022337252   0.4873704330482942   0.0018057035753268594   0.6290360757518236   0.9239031673965024   0.6030244316315164   0.8628932367593237   0.42823757101240206   0.7775185635495757   0.9175568200440535   0.6189978427050765   0.8262383748919035   0.7809858900065266   0.6510839059592866   0.032598885818912196   0.05838432027849428   0.14760475282116067   0.29985633453012367   0.552471797723999   0.9629418738819876   0.3439868761071361   0.6124876900846926   0.12452856386041002   0.80996179901957   0.39167685376988404   0.12511725703639845   0.12272286028508315   0.18092572326774636   0.4677736863733816   0.522092825404882   0.2598296235257594   0.7526881522553442   0.690255122823806   0.6045360053608285   0.6408317808206828   0.9264497773634408   0.9092692328172792   0.953452099401542   0.6082328950017707
0.8680654570849465   0.7616644799961186   0.6535957648714182   0.05576109727777161   0.9051235832029588   0.4176776038889825   0.041108074786725596   0.9312325334173616   0.09516178418338886   0.02600075011909848   0.9159908177503271   0.8085096731322784   0.9142360609156425   0.5582270637457168   0.39389799234544515   0.5486800496065191   0.1615479086602982   0.8679719409219109   0.7893619869846166   0.9078482687858361   0.23509813129685742   0.9587027081046317   0.8359098875830747   0.2996153737840655   0.3670326742119109   0.19703822810851304   0.18231412271165645   0.2438542765062939   0.461909091008952   0.7793606242195306   0.14120604792493086   0.3126217430889323   0.36674730682556317   0.753359874100432   0.2252152301746037   0.5041120699566539   0.45251124590992065   0.1951328103547152   0.8313172378291586   0.9554320203501349   0.2909633372496225   0.3271608694328043   0.04195525084454193   0.04758375156429867   0.05586520595276505   0.36845816132817266   0.20604536326146725   0.7479683777802332   0.6888325317408541   0.17141993321965965   0.02373124054981079   0.5041141012739392   0.22692344073190213   0.39205930900012914   0.8825251926248799   0.19149235818500693   0.860176133906339   0.638699434899697   0.6573099624502763   0.6873802882283531   0.4076648879964183   0.44356662454498186   0.8259927246211177   0.7319482678782182
0.11670155074679585   0.11640575511217756   0.7840374737765757   0.6843645163139195   0.0608363447940308   0.7479475937840049   0.5779921105151086   0.9363961385336863   0.37200381305317665   0.5765276605643452   0.5542608699652978   0.4322820372597471   0.1450803723212745   0.18446835156421612   0.6717356773404178   0.2407896790747402   0.2849042384149355   0.5457689166645191   0.01442571489014154   0.5534093908463872   0.8772393504185172   0.10220229211953719   0.18843299026902385   0.821461122968169   0.7605377996717214   0.9857965370073596   0.4043955164924481   0.1370966066542495   0.6997014548776905   0.23784894322335473   0.8264034059773395   0.20070046812056314   0.32769764182451394   0.6613212826590095   0.2721425360120418   0.768418430860816   0.18261726950323942   0.4768529310947934   0.600406858671624   0.5276287517860758   0.8977130310883039   0.9310840144302743   0.5859811437814825   0.9742193609396886   0.020473680669786675   0.8288817223107371   0.39754815351245865   0.15275823797151963   0.2599358809980653   0.8430851853033775   0.9931526370200106   0.015661631317270157   0.5602344261203748   0.6052362420800227   0.166749231042671   0.8149611631967071   0.2325367842958608   0.9439149594210132   0.8946066950306292   0.04654273233589102   0.04991951479262136   0.4670620283262199   0.29419983635900515   0.5189139805498152
0.15220648370431747   0.5359780138959456   0.7082186925775227   0.5446946196101266   0.13173280303453078   0.7070962915852085   0.310670539065064   0.39193638163860695   0.8717969220364655   0.864011106281831   0.3175179020450534   0.3762747503213368   0.31156249591609075   0.25877486420180823   0.1507686710023824   0.5613135871246298   0.07902571162022996   0.31485990478079495   0.2561619759717532   0.5147708547887387   0.029106196827608607   0.847797876454575   0.9619621396127481   0.9958568742389236   0.8768997131232912   0.31181986255862953   0.25374344703522544   0.45116225462879694   0.7451669100887603   0.6047235709734211   0.9430729079701614   0.05922587299019001   0.8733699880522948   0.7407124646915901   0.625555005925108   0.6829511226688533   0.5618074921362041   0.4819376004897819   0.47478633492272565   0.12163753554422349   0.48278178051597415   0.16707769570898695   0.21862435895097246   0.6068666807554848   0.4536755836883655   0.3192798192544119   0.25666221933822436   0.6110098065165612   0.5767758705650744   0.007459956695782351   0.00291877230299894   0.1598475518877643   0.831608960476314   0.40273638572236126   0.05984586433283747   0.1006216788975743   0.9582389724240191   0.6620239210307711   0.4342908584077294   0.41767055622872107   0.39643148028781505   0.18008632054098922   0.9595045234850037   0.29603302068449755
0.913649699771841   0.013008624832002257   0.7408801645340313   0.6891663399290128   0.4599741160834754   0.6937288055775904   0.4842179451958069   0.07815653341245155   0.883198245518401   0.6862688488818081   0.481299172892808   0.9183089815246872   0.051589285042086944   0.28353246315944675   0.4214533085599705   0.817687302627113   0.09335031261806777   0.6215085421286756   0.9871624501522411   0.40001674639839185   0.6969188323302528   0.4414222215876864   0.027657926667237338   0.10398372571389432   0.7832691325584118   0.42841359675568413   0.28677776213320605   0.41481738578488153   0.3232950164749364   0.7346847911780937   0.8025598169373992   0.33666085237243   0.44009677095653543   0.04841594229628573   0.3212606440445912   0.4183518708477427   0.3885074859144485   0.764883479136839   0.8998073354846207   0.6006645682206299   0.2951571732963807   0.14337493700816334   0.9126448853323796   0.20064782182223795   0.598238340966128   0.701952715420477   0.8849869586651423   0.09666409610834362   0.8149692084077163   0.2735391186647928   0.5982091965319363   0.6818467103234621   0.4916741919327798   0.538854327486699   0.7956493795945371   0.3451858579510321   0.05157742097624434   0.49043838519041333   0.4743887355499459   0.9268339871032893   0.6630699350617959   0.7255549060535743   0.5745814000653252   0.32616941888265955
0.36791276176541515   0.582179969045411   0.6619365147329456   0.12552159706042162   0.7696744207992872   0.880227253624934   0.7769495560678034   0.028857500952078   0.9547052123915709   0.6066881349601413   0.17874035953586712   0.3470107906286159   0.46303102045879113   0.06783380747344218   0.38309097994133   0.0018249326775837851   0.4114535994825468   0.5773954222830289   0.9087022443913841   0.07499094557429442   0.748383664420751   0.8518405162294546   0.33412084432605893   0.7488215266916348   0.38047090265533584   0.26966054718404353   0.6721843295931134   0.6232999296312133   0.6107964818560487   0.3894332935591095   0.89523477352531   0.5944424286791352   0.6560912694644778   0.7827451585989682   0.7164944139894429   0.24743163805051935   0.19306024900568663   0.7149113511255261   0.33340343404811285   0.24560670537293555   0.7816066495231399   0.1375159288424972   0.4247011896567287   0.17061575979864113   0.033222985102388865   0.28567541261304263   0.09058034533066976   0.42179423310700626   0.6527520824470531   0.016014865428999128   0.4183960157375564   0.7984943034757931   0.04195560059100434   0.6265815718698896   0.5231612422122465   0.2040518747966578   0.38586433112652657   0.8438364132709214   0.8066668282228036   0.9566202367461385   0.19280408212083994   0.12892506214539534   0.47326339417469077   0.7110135313732029
0.4111974325977001   0.9914091333028981   0.048562204517962046   0.5403977715745618   0.3779744474953112   0.7057337206898555   0.9579818591872923   0.11860353846755549   0.7252223650482582   0.6897188552608564   0.5395858434497358   0.32010923499176247   0.6832667644572539   0.06313728339096672   0.016424601237489393   0.11605736019510467   0.2974024333307273   0.21930087012004532   0.20975777301468582   0.1594371234489662   0.10459835120988738   0.09037580797464999   0.736494378839995   0.4484235920757633   0.6934009186121872   0.09896667467175184   0.687932174322033   0.9080258205012015   0.31542647111687605   0.39323295398189634   0.7299503151347407   0.7894222820336461   0.5902041060686178   0.70351409872104   0.1903644716850049   0.4693130470418836   0.906937341611364   0.6403768153300733   0.17393987044751552   0.35325568684677894   0.6095349082806367   0.4210759452100279   0.9641820974328297   0.1938185633978127   0.5049365570707494   0.33070013723537794   0.22768771859283463   0.7453949713220493   0.811535638458562   0.2317334625636261   0.5397555442708016   0.8373691508208478   0.496109167341686   0.8385005085817298   0.8098052291360608   0.047946868787201835   0.9059050612730681   0.13498640986068977   0.619440757451056   0.5786338217453183   0.9989677196617042   0.49460959453061654   0.4455008870035404   0.22537813489853933
0.3894328113810675   0.07353364932058862   0.4813187895707107   0.031559571500726635   0.8844962543103182   0.7428335120852106   0.2536310709778761   0.28616460017867723   0.07296061585175613   0.5111000495215846   0.7138755267070745   0.44879544935782933   0.5768514485100701   0.6725995409398549   0.9040702975710136   0.4008485805706275   0.670946387237002   0.5376131310791651   0.2846295401199577   0.8222147588253093   0.6719786675752978   0.04300353654854854   0.8391286531164173   0.59683662392677   0.28254585619423034   0.9694698872279599   0.3578098635457066   0.5652770524260433   0.3980496018839122   0.22663637514274926   0.10417879256783048   0.2791124522473661   0.3250889860321561   0.7155363256211646   0.390303265860756   0.8303170028895367   0.7482375375220859   0.0429367846813098   0.4862329682897423   0.4294684223189092   0.07729115028508395   0.5053236536021447   0.20160342816978455   0.6072536634935999   0.4053124827097861   0.4623201170535962   0.3624747750533672   0.010417039566829975   0.12276662651555575   0.49285022982563625   0.004664911507660671   0.4451399871407867   0.7247170246316436   0.266213854682887   0.9004861189398302   0.16602753489342062   0.3996280385994875   0.5506775290617224   0.5101828530790742   0.3357105320038839   0.6513905010774016   0.5077407443804126   0.023949884789331934   0.9062421096849748
0.5740993507923177   0.002417090778267834   0.8223464566195474   0.2989884461913748   0.16878686808253152   0.5400969737246717   0.45987168156618013   0.28857140662454484   0.04602024156697577   0.047246743899035396   0.45520677005851945   0.8434314194837582   0.3213032169353322   0.7810328892161483   0.5547206511186893   0.6774038845903375   0.9216751783358447   0.230355360154426   0.04453779803961502   0.34169335258645367   0.27028467725844313   0.7226146157740134   0.020587913250283092   0.4354512429014789   0.6961853264661255   0.7201975249957456   0.19824145663073572   0.13646279671010406   0.527398458383594   0.18010055127107397   0.7383697750645556   0.8478913900855592   0.4813782168166182   0.13285380737203858   0.28316300500603614   0.004459970601801028   0.16007499988128598   0.3518209181558902   0.7284423538873469   0.32705608601146346   0.2383998215454413   0.12146555800146418   0.6839045558477319   0.9853627334250098   0.9681151442869982   0.3988509422274507   0.6633166425974488   0.5499114905235309   0.27192981782087267   0.6786534172317051   0.46507518596671305   0.41344869381342686   0.7445313594372787   0.49855286596063114   0.7267054109021575   0.5655573037278676   0.26315314262066053   0.36569905858859253   0.4435424058961213   0.5610973331260666   0.10307814273937455   0.013878140432702343   0.7151000520087745   0.23404124711460314
0.8646783211939333   0.8924125824312381   0.03119549616104254   0.24867851368959332   0.8965631769069351   0.49356164020378746   0.36787885356359373   0.6987670231660624   0.6246333590860624   0.8149082229720823   0.9028036675968807   0.28531832935263557   0.8801019996487838   0.31635535701145123   0.17609825669472323   0.719761025624768   0.6169488570281232   0.9506562984228587   0.732555850798602   0.1586636924987013   0.5138707142887486   0.9367781579901563   0.017455798789827504   0.9246224453840981   0.6491923930948154   0.04436557555891816   0.986260302628785   0.6759439316945048   0.7526292161878803   0.5508039353551307   0.6183814490651912   0.9771769085284424   0.12799585710181785   0.7358957123830484   0.7155777814683105   0.6918585791758068   0.24789385745303413   0.4195403553715972   0.5394795247735873   0.972097553551039   0.630945000424911   0.4688840569487385   0.8069236739749853   0.8134338610523376   0.11707428613616229   0.5321058989585822   0.7894678751851578   0.8888114156682395   0.4678818930413469   0.48774032339966406   0.8032075725563729   0.21286748397373467   0.7152526768534666   0.9369363880445333   0.1848261234911817   0.23569057544529226   0.5872568197516488   0.20104067566148492   0.4692483420228712   0.5438319962694854   0.3393629622986146   0.7815003202898878   0.929768817249284   0.5717344427184464
0.7084179618737036   0.3126162633411492   0.12284514327429853   0.7583005816661088   0.5913436757375414   0.780510364382567   0.33337726808914064   0.8694891659978693   0.12346178269619448   0.29277004098290305   0.5301696955327677   0.6566216820241346   0.40820910584272785   0.3558336529383697   0.34534357204158606   0.42093110657884236   0.8209522860910791   0.1547929772768848   0.8760952300187149   0.8770991103093569   0.4815893237924645   0.37329265698699704   0.946326412769431   0.3053646675909105   0.7731713619187608   0.06067639364584778   0.8234812694951325   0.5470640859248017   0.18182768618121944   0.2801660292632807   0.4901040014059918   0.6775749199269324   0.058365903485024954   0.9873959882803777   0.959934305873224   0.020953237902797805   0.6501567976422971   0.631562335342008   0.614590733831638   0.6000221313239554   0.829204511551218   0.4767693580651232   0.7384955038129231   0.7229230210145985   0.3476151877587535   0.10347670107812618   0.7921690910434921   0.41755835342368797   0.5744438258399927   0.042800307432278396   0.9686878215483596   0.8704942674988863   0.39261613965877323   0.7626342781689976   0.47858382014236783   0.19291934757195378   0.33425023617374827   0.77523828988862   0.5186495142691437   0.171966109669156   0.6840934385314512   0.143675954546612   0.9040587804375059   0.5719439783452005
0.8548889269802332   0.6669065964814888   0.16556327662458276   0.8490209573306021   0.5072737392214797   0.5634298954033626   0.37339418558109067   0.43146260390691415   0.932829913381487   0.5206295879710842   0.404706364032731   0.5609683364080279   0.5402137737227138   0.7579953098020865   0.9261225438903632   0.3680489888360741   0.20596353754896554   0.9827570199134665   0.40747302962121945   0.19608287916691816   0.5218700990175144   0.8390810653668546   0.5034142491837136   0.6241389008217176   0.6669811720372811   0.17217446888536578   0.3378509725591309   0.7751179434911155   0.15970743281580144   0.6087445734820032   0.9644567869780402   0.3436553395842014   0.2268775194343144   0.08811498551091895   0.5597504229453092   0.7826870031761735   0.6866637457116006   0.33011967570883244   0.6336278790549459   0.41463801434009934   0.48070020816263503   0.34736265579536585   0.22615484943372646   0.21855513517318118   0.9588301091451207   0.5082815904285113   0.7227406002500129   0.5944162343514636   0.29184893710783955   0.33610712154314554   0.384889627690882   0.819298290860348   0.1321415042920381   0.7273625480611423   0.42043284071284176   0.47564295127614664   0.9052639848577237   0.6392475625502234   0.8606824177675326   0.6929559480999732   0.21860023914612314   0.309127886841391   0.22705453871258668   0.27831793375987385
0.7379000309834881   0.9617652310460251   0.0008996892788601949   0.05976279858669265   0.7790699218383674   0.45348364061751384   0.27815908902884734   0.4653465642352291   0.4872209847305279   0.11737651907436833   0.8932694613379654   0.646048273374881   0.3550794804384898   0.390013971013226   0.4728366206251236   0.1704053220987344   0.4498154955807661   0.7507664084630026   0.612154202857591   0.47744937399876125   0.23121525643464294   0.4416385216216116   0.38509966414500435   0.1991314402388874   0.49331522545115486   0.4798732905755865   0.38419997486614416   0.13936864165219476   0.7142453036127874   0.026389649958072643   0.10604088583729682   0.6740220774169656   0.2270243188822595   0.9090131308837043   0.21277142449933142   0.027973804042084632   0.8719448384437697   0.5189991598704783   0.7399348038742078   0.8575684819433502   0.42212934286300363   0.7682327514074757   0.12778060101661678   0.380119107944589   0.19091408642836066   0.32659422978586417   0.7426809368716124   0.1809876677057016   0.6975988609772058   0.8467209392102777   0.35848096200546825   0.04161902605350684   0.9833535573644184   0.820331289252205   0.25244007616817143   0.3675969486365412   0.7563292384821589   0.9113181583685007   0.03966865166884001   0.3396231445944565   0.8843844000383893   0.3923189984980224   0.2997338477946322   0.4820546626511063
0.4622550571753856   0.6240862470905466   0.17195324677801543   0.10193555470651731   0.27134097074702496   0.29749201730468244   0.42927230990640297   0.9209478870008158   0.5737421097698191   0.4507710780944048   0.07079134790093473   0.8793288609473089   0.5903885524054007   0.6304397888421998   0.8183512717327633   0.5117319123107678   0.8340593139232417   0.719121630473699   0.7786826200639233   0.17210876771631117   0.9496749138848525   0.32680263197567666   0.47894877226929106   0.6900541050652048   0.4874198567094669   0.7027163848851301   0.3069955254912757   0.5881185503586875   0.21607888596244196   0.4052243675804476   0.8777232155848727   0.6671706633578719   0.6423367761926229   0.9544532894860428   0.8069318676839379   0.787841802410563   0.051948223787222185   0.3240135006438431   0.9885805959511746   0.27610989009979525   0.21788890986398043   0.604891870170144   0.20989797588725134   0.1040011223834841   0.26821399597912793   0.27808923819446735   0.7309492036179602   0.4139470173182792   0.780794139269661   0.5753728533093373   0.4239536781266846   0.8258284669595917   0.5647152533072191   0.17014848572888966   0.546230462541812   0.15865780360171983   0.9223784771145962   0.21569519624284683   0.7392985948578741   0.3708160011911569   0.870430253327374   0.8916816955990038   0.7507179989066994   0.0947061110913616
0.6525413434633935   0.2867898254288597   0.5408200230194481   0.9907049887078775   0.38432734748426567   0.008700587234392387   0.8098708194014878   0.5767579713895983   0.6035332082146047   0.43332773392505514   0.38591714127480314   0.7509295044300066   0.038817954907385585   0.26317924819616545   0.8396866787329912   0.5922717008282868   0.1164394777927894   0.047484051953318646   0.10038808387511713   0.22145569963712994   0.2460092244654154   0.15580235635431489   0.3496700849684177   0.12674958854576834   0.5934678810020219   0.8690125309254552   0.8088500619489697   0.13604459983789086   0.2091405335177562   0.8603119436910628   0.9989792425474819   0.5592866284482926   0.6056073253031515   0.42698420976600765   0.6130621012726788   0.808357124018286   0.5667893703957659   0.1638049615698422   0.7733754225396876   0.21608542318999913   0.4503498926029766   0.11632090961652355   0.6729873386645704   0.9946297235528692   0.20434066813756116   0.9605185532622087   0.3233172536961527   0.8678801350071008   0.6108727871355393   0.09150602233675348   0.514467191747183   0.73183553516921   0.40173225361778314   0.2311940786456907   0.5154879491997011   0.1725489067209174   0.7961249283146316   0.804209868879683   0.9024258479270224   0.3641917827026315   0.22933555791886562   0.6404049073098408   0.12905042538733477   0.14810635951263237
0.7789856653158891   0.5240839976933173   0.45606308672276435   0.15347663595976319   0.5746449971783278   0.5635654444311087   0.13274583302661164   0.28559650095266237   0.9637722100427886   0.47205942209435514   0.6182786412794287   0.5537609657834524   0.5620399564250054   0.24086534344866445   0.10279069207972749   0.38121205906253497   0.7659150281103738   0.4366554745689814   0.20036484415270514   0.0170202763599035   0.5365794701915082   0.7962505672591406   0.07131441876537037   0.8689139168472712   0.7575938048756191   0.2721665695658233   0.6152513320426061   0.7154372808875079   0.18294880769729127   0.7086011251347146   0.4825054990159944   0.42984077993484554   0.2191765976545027   0.2365417030403595   0.8642268577365658   0.8760798141513931   0.6571366412294973   0.9956763595916951   0.7614361656568382   0.49486775508885816   0.8912216131191235   0.5590208850227136   0.5610713215041332   0.47784747872895467   0.35464214292761526   0.7627703177635731   0.48975690273876277   0.6089335618816836   0.5970483380519961   0.49060374819774977   0.8745055706961568   0.8934962809941756   0.4140995303547048   0.782002623063035   0.3920000716801623   0.46365550105933007   0.1949229327002021   0.5454609200226755   0.5277732139435966   0.5875756869079369   0.5377862914707048   0.5497845604309806   0.7663370482867583   0.09270793181907874
0.6465646783515814   0.9907636754082669   0.2052657267826251   0.614860453090124   0.29192253542396607   0.2279933576446939   0.7155088240438623   0.005926891208440565   0.69487419737197   0.7373896094469441   0.8410032533477055   0.11243061021426497   0.28077466701726517   0.9553869863839091   0.4490031816675432   0.648775109154935   0.0858517343170631   0.40992606636123347   0.9212299677239467   0.061199422246998036   0.5480654428463583   0.860141505930253   0.15489291943718844   0.9684914904279193   0.9015007644947769   0.869377830521986   0.9496271926545633   0.3536310373377952   0.6095782290708108   0.6413844728772922   0.234118368610701   0.34770414612935463   0.9147040316988408   0.903994863430348   0.3931151152629954   0.23527353591508965   0.6339293646815757   0.9486078770464389   0.9441119335954522   0.5864984267601547   0.5480776303645126   0.5386818106852055   0.02288196587150551   0.5252990045131567   0.000012187518154285195   0.6785403047549525   0.8679890464343171   0.5568075140852374   0.09851142302337733   0.8091624742329665   0.9183618537797538   0.20317647674744221   0.48893319395256646   0.16777800135567442   0.6842434851690528   0.8554723306180876   0.5742291622537257   0.2637831379253264   0.2911283699060573   0.6201987947029979   0.94029979757215   0.3151752608788875   0.3470164363106051   0.03370036794284318
0.39222216720763736   0.776493450193682   0.3241344704390996   0.5084013634296864   0.39220997968948307   0.09795314543872942   0.4561454240047825   0.9515938493444491   0.2936985566661058   0.28879067120576285   0.5377835702250288   0.7484173725970069   0.8047653627135393   0.12101266985008846   0.853540085055976   0.8929450419789193   0.23053620045981366   0.857229531924762   0.5624117151499187   0.2727462472759214   0.2902364028876637   0.5420542710458746   0.21539527883931367   0.2390458793330782   0.8980142356800264   0.7655608208521927   0.891260808400214   0.7306445159033917   0.5058042559905432   0.6676076754134632   0.4351153843954316   0.7790506665589426   0.21210569932443749   0.37881700420770037   0.8973318141704029   0.030633293961935783   0.4073403366108982   0.2578043343576119   0.0437917291144268   0.13768825198301649   0.17680413615108456   0.4005748024328498   0.481380013964508   0.8649420047070951   0.8865677332634209   0.8585205313869753   0.2659847351251944   0.625896125374017   0.9885534975833945   0.09295971053478257   0.3747239267249803   0.8952516094706252   0.48274924159285126   0.42535203512131936   0.9396085423295487   0.11620094291168252   0.27064354226841375   0.04653503091361898   0.042276728159145835   0.08556764894974674   0.8633032056575155   0.7887306965560071   0.998484999044719   0.9478793969667303
0.686499069506431   0.38815589412315726   0.517104985080211   0.08293739225963515   0.7999313362430102   0.5296353627361821   0.2511202499550166   0.45704126688561825   0.8113778386596157   0.4366756522013995   0.8763963232300364   0.5617896574149931   0.3286285970667644   0.011323617080080142   0.9367877809004876   0.44558871450331056   0.057985054798350665   0.9647885861664611   0.8945110527413418   0.3600210655535638   0.19468184914083514   0.17605788961045407   0.8960260536966228   0.41214166858683354   0.5081827796344042   0.7879019954872968   0.3789210686164118   0.3292042763271984   0.708251443391394   0.2582666327511148   0.1278008186613952   0.8721630094415802   0.8968736047317784   0.8215909805497152   0.2514044954313589   0.31037335202658706   0.568245007665014   0.8102673634696351   0.3146167145308712   0.8647846375232765   0.5102599528666633   0.845478777303174   0.4201056617895294   0.5047635719697128   0.3155781037258282   0.6694208876927199   0.5240796080929065   0.09262190338287918   0.807395324091424   0.8815188922054231   0.1451585394764948   0.7634176270556807   0.09914388070002998   0.6232522594543083   0.01735772081509958   0.8912546176141006   0.20227027596825162   0.801661278904593   0.7659532253837407   0.5808812655875135   0.6340252683032377   0.9913939154349579   0.4513365108528695   0.716096628064237
0.12376531543657435   0.1459151381317839   0.03123084906334011   0.21133305609452427   0.8081872117107461   0.476494250439064   0.5071512409704335   0.11871115271164509   0.0007918876193221843   0.5949753582336409   0.36199270149393875   0.35529352565596434   0.9016480069192923   0.9717230987793326   0.34463498067883913   0.4640389080418637   0.6993777309510406   0.17006181987473956   0.5786817552950985   0.8831576424543501   0.06535246264780295   0.17866790443978167   0.12734524444222894   0.1670610143901132   0.9415871472112286   0.032752766307997776   0.09611439537888883   0.955727958295589   0.13339993550048243   0.5562585158689338   0.5889631544084553   0.8370168055839439   0.13260804788116023   0.9612831576352929   0.2269704529145166   0.48172327992797953   0.23096004096186804   0.9895600588559603   0.8823354722356774   0.017684371886115824   0.5315823100108275   0.8194982389812208   0.303653716940579   0.13452672943176563   0.4662298473630245   0.6408303345414391   0.17630847249835008   0.9674657150416525   0.5246427001517959   0.6080775682334413   0.08019407711946125   0.011737756746063518   0.39124276465131347   0.05181905236450751   0.49123092271100594   0.17472095116211966   0.2586347167701532   0.09053589472921462   0.2642604697964894   0.6929976712341401   0.0276746758082852   0.10097583587325432   0.3819249975608119   0.6753132993480243
0.49609236579745775   0.28147759689203355   0.0782712806202329   0.5407865699162586   0.02986251843443328   0.6406472623505944   0.9019628081218828   0.5733208548746063   0.5052198182826374   0.032569694117153165   0.8217687310024215   0.5615830981285427   0.11397705363132393   0.9807506417526457   0.33053780829141566   0.386862146966423   0.8553423368611707   0.8902147470234311   0.0662773384949263   0.6938644757322829   0.8276676610528855   0.7892389111501767   0.6843523409341143   0.018551176384258582   0.3315752952554277   0.5077613142581432   0.6060810603138815   0.4777646064679999   0.30171277682099445   0.8671140519075486   0.7041182521919986   0.9044437515933937   0.7964929585383571   0.8345443577903955   0.8823495211895771   0.342860653464851   0.6825159049070332   0.8537937160377499   0.5518117128981614   0.955998506498428   0.8271735680458624   0.9635789690143188   0.48553437440323516   0.26213403076614505   0.9995059069929769   0.1743400578641421   0.8011820334691208   0.24358285438188648   0.6679306117375492   0.666578743605999   0.19510097315523925   0.7658182479138865   0.36621783491655474   0.7994646916984502   0.4909827209632406   0.8613744963204929   0.5697248763781977   0.9649203339080548   0.6086331997736635   0.5185138428556418   0.8872089714711645   0.11112661787030488   0.056821486875502085   0.562515336357214
0.060035403425302114   0.14754764885598604   0.5712871124722669   0.30038130559106885   0.06052949643232518   0.973207590991844   0.7701050790031462   0.05679845120918236   0.392598884694776   0.30662884738584495   0.575004105847907   0.2909802032952958   0.02638104977822123   0.5071641556873947   0.08402138488466633   0.4296057069748029   0.45665617340002357   0.5422438217793399   0.47538818511100284   0.911091864119161   0.569447201928859   0.4311172039090351   0.41856669823550074   0.3485765277619471   0.5094117985035569   0.283569555053049   0.8472795857632338   0.04819522217087825   0.4488823020712317   0.3103619640612051   0.0771745067600876   0.9913967709616959   0.056283417376455744   0.003733116675360125   0.5021704009121807   0.7004165676664001   0.029902367598234513   0.49656896098796544   0.4181490160275143   0.2708108606915972   0.573246194198211   0.9543251392086255   0.9427608309165115   0.35971899657243617   0.003798992269351962   0.5232079352995904   0.5241941326810108   0.011142468810489081   0.4943871937657951   0.23963838024654144   0.676914546917777   0.9629472466396108   0.04550489169456336   0.9292764161853364   0.5997400401576893   0.971550475677915   0.9892214743181076   0.9255432995099763   0.09756963924550872   0.2711339080115148   0.9593191067198731   0.4289743385220108   0.6794206232179945   0.00032304731991764286
0.38607291252166215   0.4746491993133853   0.7366597923014829   0.6406040507474815   0.38227392025231016   0.9514412640137948   0.21246565962047215   0.6294615819369924   0.8878867264865151   0.7118028837672534   0.5355511127026952   0.6665143352973816   0.8423818347919517   0.782526467581917   0.9358110725450057   0.6949638596194666   0.8531603604738441   0.8569831680719407   0.8382414332994971   0.4238299516079518   0.893841253753971   0.42800882954992997   0.15882081008150264   0.4235069042880341   0.5077683412323089   0.9533596302365447   0.42216101778001974   0.7829028535405527   0.12549442097999872   0.001918366222749854   0.2096953581595476   0.15344127160356028   0.23760769449348362   0.29011548245549645   0.6741442454568524   0.4869269363061787   0.3952258597015319   0.5075890148735794   0.7383331729118466   0.7919630766867121   0.5420654992276878   0.6506058468016387   0.9000917396123496   0.36813312507876034   0.6482242454737167   0.22259701725170866   0.741270929530847   0.9446262207907262   0.1404559042414078   0.269237387015164   0.3191099117508272   0.16172336725017358   0.014961483261409083   0.2673190207924141   0.10941455359127965   0.008282095646613297   0.7773537887679255   0.9772035383369176   0.43527030813442724   0.5213551593404345   0.3821279290663936   0.4696145234633382   0.6969371352225806   0.7293920826537225
0.8400624298387058   0.8190086766616995   0.796845395610231   0.3612589575749621   0.19183818436498914   0.596411659409991   0.055574466079384044   0.41663273678423585   0.051382280123581335   0.32717427239482694   0.7364645543285568   0.2549093695340623   0.036420796862172256   0.059855251602412854   0.6270500007372771   0.246627273887449   0.2590670080942468   0.08265171326549521   0.19177969260284994   0.7252721145470145   0.8769390790278532   0.613037189802157   0.49484255738026933   0.995880031893292   0.036876649189147355   0.7940285131404574   0.6979971617700383   0.6346210743183299   0.8450384648241582   0.19761685373046653   0.6424226956906544   0.217988337534094   0.7936561847005769   0.8704425813356396   0.9059581413620975   0.9630789680000317   0.7572353878384046   0.8105873297332267   0.27890814062482033   0.7164516941125827   0.49816837974415784   0.7279356164677315   0.08712844802197037   0.9911795795655682   0.6212293007163047   0.1148984266655745   0.592285890641701   0.9952995476722762   0.5843526515271573   0.32086991352511707   0.8942887288716627   0.3606784733539464   0.7393141867029991   0.12325305979465054   0.25186603318100836   0.1426901358198524   0.9456580020024222   0.25281047845901095   0.3459078918189109   0.1796111678198207   0.18842261416401757   0.4422231487257843   0.06699975119409057   0.46315947370723803
0.6902542344198598   0.7142875322580527   0.9798713031721202   0.47197989414166974   0.06902493370355511   0.5993891055924783   0.38758541253041917   0.47668034646939345   0.48467228217639785   0.2785191920673612   0.4932966836587565   0.11600187311544703   0.7453580954733988   0.1552661322727107   0.24143065047774814   0.9733117372955946   0.7997000934709766   0.9024556538136997   0.8955227586588372   0.7937005694757739   0.6112774793069591   0.46023250508791547   0.8285230074647467   0.3305410957685359   0.9210232448870993   0.7459449728298627   0.8486517042926265   0.8585612016268661   0.8519983111835442   0.1465558672373844   0.4610662917622073   0.3818808551574727   0.36732602900714634   0.8680366751700231   0.9677696081034508   0.26587898204202565   0.6219679335337476   0.7127705428973126   0.7263389576257027   0.29256724474643103   0.822267840062771   0.8103148890836128   0.8308161989668654   0.49886667527065715   0.21099036075581193   0.35008238399569735   0.002293191502118725   0.16832557950212124   0.2899671158687126   0.6041374111658346   0.15364148720949225   0.30976437787525507   0.4379688046851684   0.4575815439284503   0.692575195447285   0.9278835227177824   0.07064277567802205   0.589544868758427   0.7248055873438342   0.6620045406757568   0.4486748421442745   0.8767743258611146   0.9984666297181315   0.36943729592932567
0.6264070020815035   0.06645943677750177   0.16765043075126612   0.8705706206586685   0.4154166413256916   0.7163770527818044   0.16535723924914741   0.7022450411565473   0.125449525456979   0.1122396416159697   0.01171575203965515   0.3924806632812922   0.6874807207718105   0.6546580976875195   0.3191405565923702   0.4645971405635098   0.6168379450937885   0.06511322892909234   0.594334969248536   0.8025925998877531   0.16816310294951403   0.18833890306797776   0.5958683395304045   0.43315530395842744   0.5417561008680105   0.12187946629047601   0.42821790877913835   0.562584683299759   0.12633945954231893   0.4055024135086716   0.26286066952999093   0.8603396421432117   0.000889934085339951   0.2932627718927019   0.2511449174903358   0.4678589788619194   0.3134092133135294   0.6386046742051825   0.9320043608979656   0.003261838298409582   0.6965712682197408   0.5734914452760901   0.3376693916494296   0.20066923841065645   0.5284081652702268   0.38515254220811235   0.7418010521190251   0.767513934452229   0.9866520644022163   0.2632730759176363   0.31358314333988674   0.20492925115247007   0.8603126048598974   0.8577706624089647   0.05072247380989581   0.34458960900925845   0.8594226707745574   0.5645078905162628   0.79957755631956   0.876730630147339   0.546013457461028   0.9259032163110803   0.8675731954215944   0.8734687918489294
0.8494421892412871   0.3524117710349902   0.5299038037721648   0.672799553438273   0.32103402397106034   0.9672592288268779   0.7881027516531397   0.905285618986044   0.3343819595688441   0.7039861529092415   0.4745196083132529   0.7003563678335739   0.47406935470894673   0.8462154905002768   0.4237971345033571   0.35576675882431547   0.6146466839343893   0.28170759998401396   0.6242195781837971   0.4790361286769764   0.06863322647336127   0.3558043836729336   0.7566463827622028   0.605567336828047   0.21919103723207412   0.003392612637943395   0.2267425789900379   0.9327677833897741   0.8981570132610137   0.03613338381106552   0.4386398273368982   0.027482164403730053   0.5637750536921697   0.33214723090182396   0.9641202190236453   0.32712579657015617   0.08970569898322299   0.4859317404015472   0.5403230845202882   0.9713590377458406   0.4750590150488337   0.2042241404175332   0.9161035063364911   0.4923229090688642   0.4064257885754724   0.8484197567445996   0.15945712357428835   0.8867555722408172   0.1872347513433983   0.8450271441066561   0.9327145445842504   0.9539877888510432   0.2890777380823845   0.8088937602955907   0.49407471724735225   0.9265056244473131   0.7253026843902148   0.47674652939376666   0.529954498223707   0.5993798278771569   0.6355969854069918   0.9908147889922195   0.9896314137034188   0.6280207901313163
0.1605379703581582   0.7865906485746863   0.07352790736692773   0.1356978810624521   0.7541121817826858   0.9381708918300867   0.9140707837926394   0.24894230882163487   0.5668774304392875   0.09314374772343052   0.981356239208389   0.2949545199705917   0.27779969235690294   0.28424998742783986   0.4872815219610367   0.3684488955232786   0.5524970079666881   0.8075034580340732   0.9573270237373298   0.7690690676461216   0.9169000225596963   0.8166886690418537   0.967695610033911   0.14104827751480528   0.7563620522015381   0.03009802046716739   0.8941677026669832   0.0053503964523532   0.002249870418852252   0.09192712863708068   0.9800969188743439   0.7564080876307183   0.43537243997956476   0.9987833809136502   0.9987406796659549   0.46145356766012663   0.15757274762266182   0.7145333934858102   0.5114591577049182   0.09300467213684804   0.6050757396559737   0.9070299354517372   0.5541321339675884   0.32393560449072645   0.6881757170962776   0.09034126640988344   0.5864365239336775   0.18288732697592117   0.9318136648947395   0.06024324594271604   0.6922688212666942   0.17753693052356798   0.9295637944758872   0.9683161173056354   0.7121719023923504   0.42112884289284963   0.49419135449632245   0.9695327363919852   0.7134312227263955   0.959675275232723   0.33661860687366063   0.25499934290617493   0.20197206502147722   0.866670603095875
0.7315428672176869   0.3479694074544378   0.6478399310538887   0.5427349986051485   0.04336715012140938   0.25762814104455434   0.061403407120211265   0.3598476716292274   0.11155348522666991   0.19738489510183832   0.36913458585351705   0.1823107411056594   0.18198969075078267   0.22906877779620297   0.6569626834611667   0.7611818982128098   0.6877983362544602   0.25953604140421777   0.9435314607347712   0.8015066229800867   0.3511797293807996   0.00453669849804286   0.741559395713294   0.9348360198842117   0.6196368621631126   0.6565672910436051   0.09371946465940524   0.39210102127906327   0.5762697120417033   0.3989391499990507   0.03231605753919397   0.032253349649835894   0.4647162268150334   0.20155425489721238   0.663181471685677   0.8499426085441765   0.2827265360642507   0.9724854771010094   0.006218788224510287   0.08876071033136676   0.5949281998097905   0.7129494356967917   0.06268732748973907   0.28725408735128005   0.24374847042899092   0.7084127371987488   0.3211279317764451   0.3524180674670683   0.6241116082658782   0.05184544615514372   0.22740846711703985   0.9603170461880051   0.047841896224174923   0.652906296156093   0.19509240957784588   0.9280636965381691   0.5831256694091416   0.4513520412588806   0.5319109378921689   0.07812108799399263   0.3003991333448908   0.4788665641578712   0.5256921496676586   0.9893603776626259
0.7054709335351004   0.7659171284610796   0.46300482217791955   0.7021062903113459   0.4617224631061094   0.057504391262330784   0.1418768904014745   0.34968822284427753   0.8376108548402312   0.0056589451071870685   0.9144684232844347   0.3893711766562725   0.7897689586160562   0.35275264895109404   0.7193760137065888   0.46130748011810335   0.20664328920691474   0.9014006076922134   0.18746507581441985   0.38318639212411076   0.9062441558620239   0.4225340435343422   0.6617729261467612   0.3938260144614849   0.2007732223269236   0.6566169150732626   0.19876810396884162   0.691719724150139   0.7390507592208142   0.5991125238109318   0.056891213567367135   0.3420315013058615   0.901439904380583   0.5934535787037448   0.1424227902829325   0.952660324649589   0.11167094576452673   0.24070092975265073   0.4230467765763437   0.49135284453148564   0.905027656557612   0.3393003220604373   0.2355817007619239   0.10816645240737488   0.9987835006955881   0.916766278526095   0.5738087746151627   0.71434043794589   0.7980102783686644   0.26014936345283246   0.3750406706463211   0.02262071379575091   0.05895951914785026   0.6610368396419006   0.3181494570789539   0.6805892124898894   0.15751961476726725   0.06758326093815584   0.17572666679602145   0.7279288878403004   0.045848669002740525   0.8268823311855051   0.7526798902196777   0.23657604330881474
0.14082101244512854   0.48758200912506783   0.5170981894577539   0.12840959090143986   0.14203751174954046   0.5708157305989727   0.9432894148425911   0.41406915295554986   0.34402723338087604   0.31066636714614027   0.56824874419627   0.391448439159799   0.28506771423302574   0.6496295275042396   0.2500992871173161   0.7108592266699096   0.1275480994657585   0.5820462665660838   0.07437262032129469   0.9829303388296092   0.08169943046301797   0.7551639353805787   0.321692730101617   0.7463542955207945   0.9408784180178894   0.26758192625551086   0.8045945406438632   0.6179447046193546   0.7988409062683489   0.6967661956565382   0.8613051258012719   0.20387555166380475   0.45481367288747293   0.38609982851039787   0.2930563816050019   0.8124271125040058   0.1697459586544472   0.7364703010061583   0.0429570944876858   0.10156788583409618   0.04219785918868869   0.15442403444007444   0.9685844741663912   0.11863754700448696   0.9604984287256707   0.3992600990594957   0.6468917440647741   0.3722832514836925   0.01962001070778127   0.13167817280398486   0.8422972034209111   0.7543385468643379   0.2207791044394323   0.43491197714744667   0.980992077619639   0.5504629952005331   0.7659654315519594   0.04881214863704881   0.6879356960146371   0.7380358826965273   0.5962194728975122   0.31234184763089057   0.6449786015269513   0.6364679968624312
0.5540216137088235   0.15791781319081613   0.6763941273605601   0.5178304498579442   0.5935231849831528   0.7586577141313204   0.02950238329578601   0.14554719837425173   0.5739031742753715   0.6269795413273356   0.18720517987487498   0.39120865150991385   0.3531240698359392   0.19206756417988885   0.20621310225523595   0.8407456563093807   0.5871586382839799   0.14325541554284005   0.5182774062405988   0.10270977361285336   0.9909391653864676   0.8309135679119495   0.8732988047136476   0.46624177675042217   0.4369175516776442   0.6729957547211334   0.19690467735308742   0.948411326892478   0.8433943666944914   0.9143380405898129   0.1674022940573014   0.8028641285182263   0.26949119241911984   0.28735849926247736   0.9801971141824264   0.4116554770083124   0.9163671225831806   0.09529093508258853   0.7739840119271905   0.5709098206989317   0.3292084842992008   0.9520355195397485   0.2557066056865916   0.4682000470860783   0.33826931891273315   0.121121951627799   0.382407800972944   0.0019582703356561515   0.901351767235089   0.44812619690666566   0.18550312361985657   0.05354694344317817   0.05795740054059763   0.5337881563168527   0.018100829562555185   0.2506828149249519   0.7884662081214777   0.24642965705437533   0.03790371538012877   0.8390273379166395   0.8720990855382971   0.1511387219717868   0.2639197034529383   0.26811751721770777
0.5428906012390963   0.1991032024320383   0.008213097766346739   0.7999174701316294   0.20462128232636312   0.0779812508042393   0.6258052967934027   0.7979591997959733   0.3032695150912741   0.6298550538975737   0.44030217317354614   0.7444122563527951   0.24531211455067647   0.09606689758072093   0.422201343610991   0.4937294414278432   0.4568459064291987   0.8496372405263456   0.3842976282308622   0.6547021035112037   0.5847468208909016   0.6984985185545588   0.12037792477792388   0.38658458629349596   0.04185621965180534   0.49939531612252047   0.11216482701157714   0.5866671161618665   0.8372349373254422   0.4214140653182812   0.4863595302181744   0.7887079163658932   0.5339654222341681   0.7915590114207075   0.046057357044628246   0.04429566001309815   0.2886533076834917   0.6954921138399865   0.6238560134336373   0.5505662185852549   0.831807401254293   0.845854873313641   0.2395583852027751   0.8958641150740512   0.24706058036339135   0.14735635475908218   0.11918046042485121   0.5092795287805553   0.205204360711586   0.6479610386365617   0.00701563341327408   0.9226124126186886   0.36796942338614375   0.2265469733182805   0.5206561031950997   0.13390449625279544   0.8340040011519756   0.434987961897573   0.47459874615047143   0.08960883623969727   0.545350693468484   0.7394958480575864   0.8507427327168342   0.5390426176544424
0.713543292214191   0.8936409747439453   0.611184347514059   0.6431785025803911   0.4664827118507997   0.7462846199848632   0.4920038870892079   0.13389897379983592   0.2612783511392137   0.09832358134830148   0.4849882536759338   0.21128656118114722   0.8933089277530699   0.871776608030021   0.9643321504808341   0.0773820649283518   0.05930492660109429   0.436788646132448   0.48973340433036266   0.9877732286886546   0.5139542331326103   0.6972927980748617   0.6389906716135285   0.4487306110342122   0.8004109409184192   0.8036518233309162   0.027806324099469412   0.8055521084538211   0.33392822906761954   0.05736720334605308   0.5358024370102615   0.6716531346539851   0.07264987792840585   0.9590436219977516   0.05081418333432775   0.4603665734728379   0.1793409501753359   0.08726701396773062   0.08648203285349365   0.38298450854448607   0.12003602357424162   0.6504783678352827   0.596748628523131   0.39521127985583154   0.6060817904416314   0.953185569760421   0.9577579569096025   0.9464806688216194   0.805670849523212   0.14953374642950473   0.929951632810133   0.14092856036779833   0.47174262045559245   0.09216654308345167   0.39414919579987157   0.4692754257138132   0.39909274252718663   0.13312292108570006   0.3433350124655438   0.00890885224097529   0.2197517923518507   0.045855907117969434   0.25685297961205017   0.6259243436964892
0.09971576877760907   0.3953775392826868   0.6601043510889192   0.23071306384065762   0.4936339783359778   0.4421919695222658   0.7023463941793167   0.28423239501903824   0.6879631288127657   0.29265822309276107   0.7723947613691836   0.14330383465123994   0.21622050835717324   0.2004916800093094   0.378245565569312   0.6740284089374268   0.8171277658299866   0.06736875892360933   0.03491055310376822   0.6651195566964514   0.5973759734781359   0.021512851805639898   0.7780575734917181   0.03919521299996226   0.49766020470052685   0.6261353125229531   0.11795322240279893   0.8084821491593046   0.004026226364549084   0.1839433430006873   0.41560682822348227   0.5242497541402664   0.31606309755178336   0.8912851199079262   0.6432120668542987   0.38094591948902645   0.09984258919461012   0.6907934398986169   0.26496650128498667   0.7069175105515997   0.2827148233646235   0.6234246809750075   0.23005594818121847   0.04179795385514825   0.6853388498864875   0.6019118291693676   0.4519983746895004   0.002602740855185995   0.18767864518596072   0.9757765166464145   0.33404515228670145   0.19412059169588136   0.18365241882141164   0.7918331736457273   0.9184383240632192   0.6698708375556149   0.8675893212696283   0.900548053737801   0.27522625720892047   0.28892491806658854   0.7677467320750182   0.20975461383918417   0.010259755923933795   0.5820074075149888
0.48503190871039464   0.5863299328641767   0.7802038077427154   0.5402094536598406   0.7996930588239071   0.9844181036948091   0.3282054330532149   0.5376067128046546   0.6120144136379464   0.00864158704839459   0.9941602807665134   0.34348612110877325   0.42836199481653475   0.21680841340266738   0.07572195670329426   0.6736152835531583   0.5607726735469064   0.3162603596648664   0.8004956994943738   0.3846903654865697   0.7930259414718883   0.1065057458256822   0.79023594357044   0.8026829579715808   0.3079940327614936   0.5201758129615055   0.01003213582772466   0.26247350431174027   0.5083009739375866   0.5357577092666964   0.6818267027745097   0.7248667915070857   0.8962865602996402   0.5271161222183018   0.6876664220079962   0.3813806703983124   0.46792456548310546   0.31030770881563446   0.611944465304702   0.7077653868451542   0.9071518919361989   0.9940473491507681   0.8114487658103282   0.32307502135858446   0.11412595046431068   0.8875416033250859   0.021212822239888234   0.5203920633870036   0.806131917702817   0.36736579036358036   0.011180686412163573   0.2579185590752634   0.2978309437652305   0.8316080810968839   0.32935398363765384   0.5330517675681777   0.4015443834655903   0.3044919588785821   0.6416875616296576   0.15167109716986532   0.9336198179824848   0.9941842500629476   0.029743096324955573   0.44390571032471116
0.02646792604628589   0.0001369009121795178   0.21829433051462735   0.12083068896612666   0.9123419755819752   0.11259529758709363   0.1970815082747391   0.600438625579123   0.10621005787915817   0.7452295072235132   0.18590082186257556   0.34252006650385963   0.8083791141139277   0.9136214261266293   0.8565468382249217   0.8094682989356818   0.40683473064833736   0.6091294672480473   0.21485927659526413   0.6577972017658166   0.47321491266585247   0.6149452171850996   0.18511618027030854   0.21389149144110542   0.4467469866195666   0.6148083162729201   0.9668218497556812   0.09306080247497878   0.5344050110375914   0.5022130186858265   0.7697403414809421   0.49262217689585575   0.4281949531584332   0.7569835114623132   0.5838395196183666   0.1501021103919961   0.6198158390445055   0.8433620853356839   0.7272926813934448   0.3406338114563142   0.21298110839616816   0.23423261808763662   0.5124334047981807   0.6828366096904976   0.7397661957303157   0.619287400902537   0.32731722452787215   0.4689451182493922   0.2930192091107491   0.004479084629616851   0.36049537477219096   0.37588431577441345   0.7586141980731577   0.5022660659437903   0.5907550332912489   0.8832621388785576   0.33041924491472446   0.7452825544814772   0.006915513672882331   0.7331600284865616   0.710603405870219   0.9019204691457933   0.2796228322794375   0.3925262170302473
0.4976222974740508   0.6676878510581566   0.7671894274812568   0.7096896073397497   0.7578561017437351   0.048400450155619626   0.43987220295338464   0.24074448909035745   0.46483689263298605   0.04392136552600278   0.07937682818119371   0.864860173315944   0.7062226945598283   0.5416552995822125   0.48862179488994484   0.9815980344373864   0.37580344964510387   0.7963727451007353   0.4817062812170625   0.24843800595082474   0.665200043774885   0.894452275954942   0.202083448937625   0.8559117889205774   0.16757774630083416   0.22676442489678544   0.4348940214563682   0.14622218158082773   0.4097216445570991   0.17836397474116583   0.9950218185029835   0.9054776924904703   0.944884751924113   0.13444260921516304   0.9156449903217898   0.04061751917452627   0.23866205736428464   0.5927873096329507   0.427023195431845   0.05901948473713997   0.8628586077191808   0.7964145645322154   0.9453169142147825   0.8105814787863153   0.19765856394429582   0.9019622885772732   0.7432334652771575   0.9546696898657379   0.030080817643461637   0.6751978636804878   0.30833944382078926   0.8084475082849101   0.6203591730863626   0.49683388893932195   0.3133176253178057   0.9029698157944398   0.6754744211622495   0.3623912797241589   0.39767263499601585   0.8623522966199135   0.4368123637979649   0.7696039700912083   0.9706494395641708   0.8033328118827736
0.5739537560787842   0.973189405558993   0.02533252534938837   0.9927513330964584   0.37629519213448837   0.07122711698171973   0.2820990600722309   0.038081643230720524   0.3462143744910267   0.3960292533012319   0.9737596162514416   0.22963413494581042   0.7258552014046641   0.8991953643619099   0.6604419909336359   0.32666431915137056   0.05038078024241457   0.536804084637751   0.2627693559376201   0.46431202253145704   0.6135684164444497   0.7672001145465427   0.2921199163734492   0.6609792106486834   0.0396146603656655   0.7940107089875497   0.26678739102406085   0.668227877552225   0.6633194682311772   0.72278359200583   0.98468833095183   0.6301462343215045   0.31710509374015045   0.3267543387045981   0.010928714700388305   0.4005120993756941   0.5912498923354863   0.42755897434268814   0.3504867237667524   0.07384778022432353   0.5408691120930718   0.8907548897049371   0.08771736782913232   0.6095357576928665   0.927300695648622   0.12355477515839444   0.7955974514556832   0.9485565470441831   0.8876860352829565   0.3295440661708447   0.5288100604316223   0.28032866949195806   0.22436656705177943   0.6067604741650148   0.5441217294797923   0.6501824351704535   0.907261473311629   0.28000613546041664   0.5331930147794041   0.24967033579475942   0.3160115809761427   0.8524471611177286   0.18270629101265168   0.17582255557043588
0.7751424688830709   0.9616922714127913   0.09498892318351934   0.5662867978775694   0.8478417732344489   0.8381374962543969   0.2993914717278362   0.6177302508333863   0.9601557379514922   0.5085934300835522   0.7705814112962139   0.33740158134142817   0.7357891708997129   0.9018329559185375   0.22645968181642157   0.6872191461709747   0.8285276975880839   0.6218268204581209   0.6932666670370174   0.43754881037621524   0.5125161166119412   0.7693796593403923   0.5105603760243659   0.2617262548057793   0.7373736477288703   0.807687387927601   0.4155714528408465   0.69543945692821   0.8895318744944214   0.969549891673204   0.11617998111301027   0.07770920609482374   0.929376136542929   0.4609564615896518   0.3455985698167964   0.7403076247533955   0.19358696564321623   0.5591235056711144   0.1191388880003748   0.05308847858242088   0.3650592680551324   0.9372966852129936   0.4258722209633573   0.6155396682062056   0.8525431514431913   0.1679170258726012   0.9153118449389914   0.35381341340042627   0.11516950371432104   0.36022963794500024   0.49974039209814497   0.6583739564722163   0.2256376292198997   0.3906797462717962   0.3835604109851347   0.5806647503773926   0.2962614926769706   0.9297232846821444   0.03796184116833835   0.840357125623997   0.10267452703375436   0.37059977901103003   0.9188229531679636   0.7872686470415762
0.737615258978622   0.4333030937980365   0.4929507322046063   0.17172897883537053   0.8850721075354308   0.2653860679254353   0.5776388872656149   0.8179155654349443   0.7699026038211096   0.905156429980435   0.07789849516746983   0.15954160896272793   0.54426497460121   0.5144766837086387   0.6943380841823351   0.5788768585853353   0.2480034819242394   0.5847533990264944   0.6563762430139968   0.7385197329613383   0.14532895489048503   0.2141536200154644   0.7375532898460332   0.9512510859197622   0.40771369591186307   0.7808505262174279   0.24460255764142694   0.7795221070843916   0.5226415883764324   0.5154644582919926   0.6669636703758122   0.9616065416494474   0.7527389845553226   0.6103080283115576   0.5890651752083423   0.8020649326867194   0.20847400995411264   0.09583134460291882   0.8947270910260071   0.2231880741013841   0.9604705280298732   0.5110779455764244   0.2383508480120104   0.4846683411400458   0.8151415731393882   0.29692432556096   0.5007975581659772   0.5334172552202837   0.40742787722752516   0.516073799343532   0.25619500052455024   0.7538951481358921   0.8847862888510928   0.0006093410515394418   0.5892313301487381   0.7922886064864447   0.13204730429577016   0.3903013127399818   0.00016615494039582865   0.9902236737997253   0.9235732943416576   0.294469968137063   0.10543906391438866   0.7670355996983411
0.9631027663117843   0.7833920225606386   0.8670882159023783   0.28236725855829536   0.1479611931723961   0.4864676969996786   0.36629065773640107   0.7489500033380116   0.7405333159448709   0.9703938976561465   0.11009565721185083   0.9950548552021196   0.8557470270937781   0.969784556604607   0.5208643270631127   0.20276624871567492   0.723699722798008   0.5794832438646252   0.5206981721227169   0.21254257491594963   0.8001264284563504   0.28501327572756224   0.41525910820832823   0.4455069752176085   0.8370236621445661   0.5016212531669236   0.54817089230595   0.16313971665931315   0.68906246897217   0.015153556167245055   0.18188023456954888   0.41418971332130144   0.9485291530272991   0.04475965851109854   0.07178457735769805   0.41913485811918183   0.09278212593352096   0.07497510190649147   0.5509202502945854   0.21636860940350694   0.369082403135513   0.4954918580418662   0.03022207817186848   0.0038260344875573017   0.5689559746791625   0.21047858231430394   0.6149629699635403   0.5583190592699488   0.7319323125345963   0.7088573291473803   0.06679207765759032   0.39517934261063564   0.04286984356242631   0.6937037729801352   0.8849118430880415   0.9809896292893342   0.0943406905351272   0.6489441144690367   0.8131272657303434   0.5618547711701524   0.0015585646016062448   0.5739690125625453   0.26220701543575803   0.3454861617666454
0.6324761614660933   0.07847715452067903   0.23198493726388958   0.3416601272790881   0.06352018678693075   0.8679985722063751   0.6170219673003493   0.7833410680091393   0.3315878742523344   0.15914124305899477   0.550229889642759   0.38816172539850363   0.2887180306899081   0.46543747007885955   0.6653180465547175   0.40717209610916943   0.19437734015478086   0.8164933556098228   0.8521907808243742   0.845317324939017   0.19281877555317462   0.2425243430472776   0.5899837653886161   0.49983116317237164   0.5603426140870813   0.16404718852659855   0.3579988281247265   0.15817103589328355   0.4968224273001506   0.2960486163202235   0.7409768608243772   0.37482996788414424   0.16523455304781623   0.1369073732612287   0.1907469711816182   0.9866682424856407   0.8765165223579081   0.6714699031823692   0.5254289246269007   0.5794961463764712   0.6821391822031273   0.8549765475725464   0.6732381438025266   0.7341788214374542   0.4893204066499527   0.6124522045252687   0.0832543784139105   0.2343476582650825   0.9289777925628714   0.44840501599867016   0.725255550289184   0.07617662237179894   0.43215536526272075   0.1523563996784467   0.9842786894648068   0.7013466544876547   0.2669208122149045   0.015449026417217992   0.7935317182831886   0.7146784120020141   0.3904042898569963   0.3439791232348488   0.2681027936562879   0.1351822656255428
0.7082651076538691   0.4890025756623025   0.5948646498537614   0.40100344418808864   0.21894470100391636   0.8765503711370338   0.5116102714398509   0.16665578592300617   0.289966908441045   0.4281453551383636   0.7863547211506668   0.09047916355120722   0.8578115431783243   0.2757889554599169   0.8020760316858601   0.3891325090635525   0.5908907309634197   0.2603399290426989   0.008544313402671444   0.6744540970615385   0.2004864411064234   0.9163608058078501   0.7404415197463835   0.5392718314359957   0.49222133345255437   0.4273582301455476   0.1455768698926221   0.13826838724790702   0.273276632448638   0.5508078590085138   0.6339665984527713   0.9716126013249009   0.983309724007593   0.12266250387015021   0.8476118773021043   0.8811334377736937   0.12549818082926872   0.8468735484102333   0.04553584561624427   0.4920009287101411   0.534607449865849   0.5865336193675343   0.03699153221357283   0.8175468316486026   0.3341210087594256   0.6701728135596843   0.2965500124671893   0.2782750002126069   0.8418996753068713   0.24281458341413673   0.1509731425745672   0.1400066129646999   0.5686230428582332   0.6920067244056229   0.517006544121796   0.16839401163979906   0.5853133188506402   0.5693442205354727   0.6693946668196916   0.28726057386610543   0.4598151380213715   0.7224706721252394   0.6238588212034474   0.7952596451559644
0.9252076881555225   0.135937052757705   0.5868672889898745   0.9777128135073617   0.5910866793960969   0.46576423919802074   0.29031727652268524   0.6994378132947549   0.7491870040892257   0.222949655783884   0.139344133948118   0.5594312003300549   0.18056396123099244   0.5309429313782611   0.622337589826322   0.39103718869025583   0.5952506423803522   0.9615987108427884   0.9529429230066304   0.10377661482415039   0.13543550435898075   0.239128038717549   0.329084101803183   0.30851696966818604   0.21022781620345823   0.103190985959844   0.7422168128133084   0.3308041561608243   0.6191411368073614   0.6374267467618233   0.45189953629062324   0.6313663428660695   0.8699541327181356   0.4144770909779393   0.31255540234250523   0.07193514253601463   0.6893901714871432   0.8835341595996782   0.6902178125161832   0.6808979538457588   0.09413952910679098   0.9219354487568897   0.7372748895095528   0.5771213390216084   0.9587040247478102   0.6828074100393408   0.4081907877063698   0.26860436935342236   0.748476208544352   0.5796164240794968   0.6659739748930613   0.937800213192598   0.1293350717369907   0.9421896773176734   0.2140744386024381   0.3064338703265285   0.259380939018855   0.5277125863397342   0.9015190362599329   0.2344987277905139   0.5699907675317119   0.644178426740056   0.21130122374374974   0.553600773944755
0.47585123842492083   0.7222429779831663   0.47402633423419693   0.9764794349231467   0.5171472136771106   0.03943556794382556   0.06583554652782715   0.7078750655697243   0.7686710051327585   0.4598191438643288   0.3998615716347658   0.7700748523771263   0.6393359333957679   0.5176294665466554   0.1857871330323277   0.4636409820505977   0.3799549943769129   0.9899168802069211   0.2842680967723948   0.22914225426008386   0.8099642268452011   0.34573845346686516   0.07296687302864505   0.6755414803153288   0.33411298842028025   0.6234954754836989   0.5989405387944481   0.6990620453921821   0.8169657747431697   0.5840599075398734   0.533104992266621   0.9911869798224578   0.04829476961041104   0.1242407636755445   0.13324342063185515   0.22111212744533154   0.40895883621464313   0.6066112971288892   0.9474562875995275   0.7574711453947338   0.029003841837730214   0.6166944169219679   0.6631881908271327   0.52832889113465   0.21903961499252914   0.27095596345510276   0.5902213177984876   0.8527874108193212   0.8849266265722489   0.6474604879714039   0.9912807790040395   0.15372536542713905   0.06796085182907925   0.06340058043153057   0.45817578673741854   0.16253838560468126   0.019666082218668206   0.939159816755986   0.3249323661055634   0.9414262581593498   0.610707246004025   0.332548519627097   0.37747607850603593   0.18395511276461593
0.5817034041662948   0.7158541027051291   0.7142878876789033   0.655626221629966   0.36266378917376574   0.44489813925002625   0.1240665698804156   0.8028388108106448   0.47773716260151683   0.7974376512786223   0.13278579087637607   0.6491134453835058   0.4097763107724376   0.7340370708470918   0.6746100041389576   0.48657505977882454   0.3901102285537694   0.7948772540911057   0.34967763803339413   0.5451488016194748   0.7794029825497443   0.46232873446400874   0.9722015595273582   0.36119368885485886   0.19769957838344943   0.7464746317588797   0.25791367184845493   0.7055674672248928   0.8350357892096837   0.3015764925088535   0.13384710196803934   0.902728656414248   0.35729862660816686   0.5041388412302311   0.0010613110916632685   0.2536152110307422   0.9475223158357292   0.7701017703831393   0.32645130695270574   0.7670401512519177   0.5574120872819598   0.9752245162920337   0.9767736689193116   0.22189134963244292   0.7780091047322155   0.5128957818280249   0.004572109391953455   0.860697660777584   0.5803095263487661   0.7664211500691452   0.7466584375434985   0.15513019355269125   0.7452737371390824   0.46484465756029175   0.6128113355754592   0.25240153713844327   0.38797511053091555   0.9607058163300606   0.6117500244837959   0.998786326107701   0.44045279469518633   0.19060404594692126   0.28529871753109015   0.23174617485578333
0.8830407074132265   0.2153795296548876   0.3085250486117785   0.009854825223340413   0.10503160268101094   0.7024837478268626   0.303952939219825   0.14915716444575633   0.5247220763322449   0.9360625977577175   0.5572945016763265   0.9940269708930651   0.7794483391931625   0.47121794019742574   0.9444831661008674   0.7416254337546219   0.3914732286622469   0.5105121238673651   0.33273314161707146   0.7428391076469208   0.9510204339670606   0.3199080779204439   0.04743442408598133   0.5110929327911374   0.06797972655383407   0.10452854826555631   0.7389093754742029   0.5012381075677971   0.9629481238728231   0.4020448004386936   0.4349564362543778   0.35208094312204075   0.4382260475405783   0.4659822026809761   0.8776619345780512   0.3580539722289756   0.6587777083474159   0.9947642624835504   0.9331787684771838   0.6164285384743537   0.26730447968516896   0.48425213861618527   0.6004456268601124   0.873589430827433   0.3162840457181084   0.16434406069574134   0.5530112027741311   0.3624964980362955   0.24830431916427437   0.059815512430185035   0.8141018272999282   0.8612583904684984   0.28535619529145123   0.6577707119914914   0.37914539104555045   0.5091774473464576   0.8471301477508729   0.19178850931051525   0.5014834564674993   0.15112347511748206   0.18835243940345708   0.19702424682696487   0.5683046879903154   0.5346949366431283
0.9210479597182881   0.7127721082107796   0.9678590611302029   0.6611055058156953   0.6047639140001797   0.5484280475150383   0.4148478583560719   0.2986090077793998   0.35645959483590534   0.48861253508485325   0.6007460310561437   0.43735061731090136   0.0711033995444541   0.8308418230933619   0.2216006400105932   0.9281731699644437   0.22397325179358116   0.6390533137828466   0.720117183543094   0.7770496948469616   0.03562081239012407   0.44202906695588173   0.15181249555277862   0.24235475820383334   0.11457285267183595   0.7292569587451021   0.18395343442257564   0.5812492523881381   0.5098089386716562   0.1808289112300638   0.7691055760665038   0.28264024460873827   0.1533493438357509   0.6922163761452106   0.16835954501036007   0.845289627297837   0.08224594429129682   0.8613745530518487   0.9467589049997669   0.9171164573333933   0.8582726924977157   0.22232123926900213   0.22664172145667288   0.14006676248643166   0.8226518801075916   0.7802921723131204   0.07482922590389428   0.8977120042825983   0.7080790274357557   0.051035213568018344   0.8908757914813187   0.31646275189446027   0.19827008876409938   0.8702063023379546   0.12177021541481489   0.033822507285722024   0.04492074492834847   0.17798992619274398   0.9534106704044548   0.18853287998788512   0.9626748006370517   0.3166153731408953   0.006651765404687952   0.27141642265449184
0.104402108139336   0.09429413387189312   0.7800100439480151   0.13134966016806018   0.2817502280317444   0.3140019615587727   0.7051808180441208   0.23363765588546187   0.5736712005959888   0.26296674799075437   0.8143050265628021   0.9171749039910015   0.37540111183188934   0.39276044565279983   0.6925348111479872   0.8833523967052795   0.3304803669035409   0.21477051946005582   0.7391241407435324   0.6948195167173944   0.36780556626648925   0.8981551463191606   0.7324723753388445   0.42340309406290255   0.26340345812715327   0.8038610124472675   0.9524623313908294   0.2920534338948424   0.9816532300954088   0.48985905088849474   0.24728151334670864   0.05841577800938051   0.4079820294994201   0.2268923028977404   0.4329764867839065   0.14124087401837893   0.03258091766753072   0.8341318572449407   0.7404416756359192   0.2578884773130994   0.7021005507639898   0.6193613377848848   0.0013175348923868493   0.563068960595705   0.3342949844975006   0.7212061914657242   0.2688451595535424   0.13966586653280236   0.07089152637034735   0.9173451790184568   0.31638282816271296   0.8476124326379599   0.0892382962749385   0.42748612812996206   0.06910131481600436   0.7891966546285795   0.6812562667755184   0.20059382523222163   0.6361248280320979   0.6479557806102005   0.6486753491079877   0.36646196798728103   0.8956831523961786   0.39006730329710115
0.9465747983439978   0.7471006302023963   0.8943656175037917   0.8269983427013962   0.6122798138464973   0.025894438736672035   0.6255204579502494   0.6873324761685938   0.54138828747615   0.10854925971821525   0.3091376297875364   0.8397200435306339   0.4521499912012114   0.6810631315882532   0.24003631497153202   0.05052338890205437   0.770893724425693   0.4804693063560316   0.6039114869394342   0.40256760829185384   0.12221837531770532   0.11400733836875053   0.7082283345432555   0.012500304994752683   0.17564357697370744   0.3669067081663543   0.8138627170394638   0.18550196229335647   0.5633637631272101   0.34101226942968227   0.18834225908921445   0.49816948612476264   0.021975475651060245   0.232463009711467   0.8792046293016781   0.6584494425941287   0.5698254844498488   0.5513998781232138   0.6391683143301461   0.6079260536920744   0.7989317600241558   0.07093057176718222   0.03525682739071191   0.20535844540022058   0.6767133847064505   0.9569232333984317   0.32702849284745633   0.1928581404054679   0.501069807732743   0.5900165252320774   0.5131657758079925   0.007356178112111422   0.9377060446055329   0.24900425580239516   0.32482351671877807   0.5091866919873488   0.9157305689544726   0.016541246090928167   0.4456188874171   0.8507372493932199   0.3459050845046238   0.4651413679677144   0.8064505730869539   0.24281119570114557
0.546973324480468   0.3942107962005322   0.771193745696242   0.03745275030092498   0.8702599397740175   0.43728756280210046   0.44416525284878566   0.8445946098954571   0.3691901320412745   0.8472710375700231   0.9309994770407931   0.8372384317833457   0.4314840874357416   0.5982667817676279   0.606175960322015   0.3280517397959969   0.515753518481269   0.5817255356766997   0.16055707290491505   0.4773144904027769   0.1698484339766452   0.11658416770898535   0.35410649981796116   0.23450329470163134   0.6228751094961772   0.7223733715084532   0.5829127541217192   0.19705054440070635   0.7526151697221597   0.28508580870635275   0.13874750127293348   0.35245593450524926   0.38342503768088526   0.43781477113632966   0.20774802423214034   0.5152175027219036   0.9519409502451437   0.8395479893687018   0.6015720639101253   0.18716576292590675   0.43618743176387464   0.2578224536920021   0.44101499100521024   0.7098512725231299   0.2663389977872294   0.14123828598301671   0.08690849118724911   0.4753479778214985   0.6434638882910522   0.41886491447456353   0.50399573706553   0.27829743342079216   0.8908487185688925   0.13377910576821078   0.3652482357925965   0.9258414989155429   0.5074236808880073   0.6959643346318811   0.15750021156045618   0.4106239961936393   0.5554827306428636   0.8564163452631793   0.5559281476503308   0.22345823326773254
0.11929529887898895   0.5985938915711773   0.11491315664512061   0.5136069607446027   0.8529563010917596   0.4573556055881605   0.028004665457871503   0.038258982923104166   0.20949241280070735   0.038490691113597014   0.5240089283923415   0.759961549502312   0.3186436942318149   0.9047115853453862   0.158760692599745   0.8341200505867691   0.8112200133438077   0.20874725071350514   0.0012604810392888304   0.42349605439312976   0.2557372827009441   0.3523309054503258   0.44533233338895795   0.20003782112539722   0.13644198382195513   0.7537370138791486   0.33041917674383736   0.6864308603807946   0.2834856827301956   0.296381408290988   0.30241451128596586   0.6481718774576903   0.07399326992948826   0.25789071717739104   0.7784055828936244   0.8882103279553784   0.7553495756976734   0.3531791318320048   0.6196448902938794   0.054090277368609316   0.9441295623538657   0.14443188111849967   0.6183844092545905   0.6305942229754795   0.6883922796529216   0.7921009756681738   0.17305207586563254   0.4305564018500823   0.5519502958309666   0.03836396178902526   0.8426328991217952   0.7441255414692878   0.2684646131007709   0.7419825534980372   0.5402183878358293   0.0959536640115974   0.19447134317128265   0.4840918363206462   0.761812804942205   0.207743336056219   0.43912176747360926   0.13091270448864137   0.14216791464832568   0.15365305868760967
0.4949922051197435   0.9864808233701418   0.5237835053937352   0.5230588357121302   0.8065999254668219   0.19437984770196787   0.35073142952810266   0.09250243386204783   0.25464962963585536   0.1560158859129426   0.5080985304063075   0.3483768923927601   0.9861850165350844   0.4140333324149054   0.9678801425704782   0.25242322838116266   0.7917136733638018   0.9299414960942592   0.20606733762827312   0.04467989232494368   0.3525919058901925   0.7990287916056178   0.06389942297994743   0.891026833637334   0.857599700770449   0.8125479682354761   0.5401159175862122   0.36796799792520385   0.0509997753036271   0.6181681205335082   0.1893844880581096   0.27546556406315603   0.7963501456677717   0.46215223462056565   0.6812859576518021   0.927088671670396   0.8101651291326873   0.04811890220566025   0.7134058150813241   0.6746654432892333   0.01845145576888553   0.11817740611140103   0.5073384774530509   0.6299855509642897   0.665859549878693   0.3191486145057832   0.4434390544731035   0.7389587173269556   0.808259849108244   0.506600646270307   0.9033231368868913   0.37099071940175177   0.7572600738046169   0.8884325257367988   0.7139386488287817   0.09552515533859572   0.9609099281368452   0.4262802911162331   0.03265269117697951   0.16843648366819977   0.15074479900415788   0.3781613889105729   0.3192468760956555   0.49377104037896646
0.13229334323527234   0.25998398279917184   0.8119083986426046   0.8637854894146769   0.4664337933565793   0.9408353682933887   0.3684693441695011   0.12482677208772129   0.6581739442483353   0.4342347220230816   0.46514620728260986   0.7538360526859695   0.9009138704437184   0.5458021962862829   0.7512075584538283   0.6583108973473738   0.9400039423068731   0.11952190517004972   0.7185548672768487   0.48987441367917406   0.7892591433027153   0.7413605162594769   0.3993079911811932   0.9961033733002076   0.656965800067443   0.481376533460305   0.5873995925385886   0.1323178838855307   0.1905320067108636   0.5405411651669163   0.2189302483690875   0.0074911117978094   0.5323580624625283   0.10630644314383471   0.7537840410864777   0.25365505911183983   0.63144419201881   0.5605042468575518   0.0025764826326494187   0.595344161764466   0.6914402497119368   0.4409823416875021   0.2840216153558007   0.10546974808529196   0.9021811064092216   0.6996218254280253   0.8847136241746075   0.10936637478508439   0.2452153063417786   0.21824529196772027   0.2973140316360189   0.9770484908995537   0.054683299630914985   0.6777041268008039   0.07838378326693138   0.9695573791017443   0.5223252371683866   0.5713976836569693   0.32459974218045373   0.7159023199899044   0.8908810451495767   0.010893436799417398   0.3220232595478043   0.12055815822543842
0.1994407954376399   0.5699110951119153   0.0380016441920036   0.015088410140146455   0.2972596890284184   0.87028926968389   0.1532880200173961   0.9057220353550621   0.05204438268663981   0.6520439777161697   0.8559739883813772   0.9286735444555084   0.9973610830557248   0.9743398509153658   0.7775902051144459   0.9591161653537641   0.47503584588733816   0.4029421672583965   0.4529904629339921   0.24321384536385965   0.5841548007377614   0.3920487304589791   0.1309672033861878   0.12265568713842123   0.3847140053001215   0.8221376353470639   0.0929655591941842   0.10756727699827479   0.08745431627170312   0.9518483656631739   0.9396775391767881   0.20184524164321271   0.03540993358506332   0.29980438794700415   0.08370355079541088   0.27317169718770434   0.0380488505293385   0.3254645370316384   0.30611334568096504   0.31405553183394025   0.5630130046420003   0.9225223697732419   0.8531228827469729   0.07084168647008059   0.9788582039042389   0.5304736393142628   0.7221556793607851   0.9481859993316594   0.5941441986041174   0.708336003967199   0.6291901201666009   0.8406187223333845   0.5066898823324143   0.7564876383040251   0.6895125809898128   0.6387734806901719   0.47127994874735096   0.45668325035702095   0.6058090301944019   0.3656017835024675   0.4332310982180124   0.13121871332538257   0.2996956845134369   0.051546251668527304
0.8702180935760121   0.20869634355214067   0.446572801766464   0.9807045651984467   0.8913598896717732   0.6782227042378779   0.7244171224056789   0.032518565866787356   0.2972156910676558   0.9698867002706789   0.09522700223907798   0.19189984353340278   0.7905258087352416   0.2133990619666538   0.40571442124926516   0.5531263628432309   0.3192458599878906   0.7567158116096329   0.7999053910548632   0.18752457934076336   0.8860147617698781   0.6254970982842503   0.5002097065414263   0.13597832767223605   0.01579666819386606   0.4168007547321096   0.05363690477496225   0.15527376247378935   0.12443677852209287   0.7385780504942316   0.32921978236928334   0.12275519660700199   0.8272210874544371   0.7686913502235527   0.23399278013020539   0.9308553530735992   0.03669527871919553   0.5552922882568989   0.8282783588809403   0.3777289902303683   0.717449418731305   0.798576476647266   0.028372967826077018   0.19020441088960494   0.8314346569614268   0.1730793783630158   0.5281632612846507   0.05422608321736889   0.8156379887675607   0.7562786236309063   0.4745263565096885   0.8989523207435796   0.6912012102454679   0.017700573136674513   0.14530657414040515   0.7761971241365776   0.8639801227910308   0.24900922291312175   0.9113137940101997   0.8453417710629784   0.8272848440718352   0.6937169346562229   0.08303543512925955   0.46761278083261004
0.10983542534053031   0.8951404580089567   0.05466246730318253   0.2774083699430051   0.27840076837910355   0.7220610796459409   0.5264992060185317   0.2231822867256362   0.46276277961154283   0.9657824560150348   0.05197284950884329   0.32422996598205667   0.771561569366075   0.9480818828783603   0.9066662753684381   0.5480328418454791   0.9075814465750442   0.6990726599652385   0.9953524813582384   0.7026910707825007   0.08029660250320896   0.005355725309015649   0.9123170462289788   0.23507828994989072   0.9704611771626787   0.11021526730005891   0.8576545789257963   0.9576699200068857   0.6920604087835751   0.38815418765411797   0.33115537290726454   0.7344876332812494   0.22929762917203225   0.42237173163908326   0.27918252339842126   0.4102576672991928   0.4577360598059573   0.474289848760723   0.37251624802998307   0.8622248254537137   0.5501546132309131   0.7752171887954845   0.3771637666717447   0.15953375467121295   0.4698580107277041   0.7698614634864689   0.46484672044276587   0.9244554647213222   0.4993968335650255   0.65964619618641   0.6071921415169695   0.9667855447144366   0.8073364247814504   0.271492008532292   0.27603676860970505   0.23229791143318718   0.5780387956094182   0.8491202768932088   0.9968542452112839   0.8220402441339943   0.12030273580346085   0.3748304281324858   0.6243379971813008   0.9598154186802808
0.5701481225725478   0.5996132393370013   0.24717423050955603   0.8002816640090678   0.10029011184484364   0.8297517758505323   0.7823275100667901   0.8758261992877455   0.6008932782798182   0.17010557966412235   0.1751353685498206   0.909040654573309   0.7935568534983678   0.8986135711318303   0.8990985999401155   0.6767427431401217   0.21551805788894962   0.04949329423862154   0.9022443547288317   0.8547024990061274   0.09521532208548879   0.6746628661061358   0.27790635754753096   0.8948870803258466   0.525067199512941   0.07504962676913454   0.030732127037974923   0.09460541631677889   0.42477708766809735   0.2452978509186022   0.24840461697118477   0.21877921702903336   0.8238838093882792   0.07519227125447987   0.07326924842136419   0.3097385624557244   0.030326955889911463   0.17657870012264956   0.17417064848124866   0.6329958193156027   0.8148088980009618   0.127085405884028   0.27192629375241695   0.7782933203094753   0.719593575915473   0.45242253977789226   0.994019936204886   0.8834062399836285   0.194526376402532   0.3773729130087577   0.963287809166911   0.7888008236668497   0.7697492887344346   0.1320750620901555   0.7148831921957263   0.5700216066378163   0.9458654793461554   0.056882790835675615   0.6416139437743621   0.26028304418209197   0.915538523456244   0.8803040907130261   0.46744329529311346   0.6272872248664894
0.10072962545528212   0.753218684828998   0.1955170015406965   0.8489939045570141   0.38113604953980906   0.3007961450511058   0.20149706533581052   0.9655876645733854   0.18660967313727705   0.9234232320423481   0.23820925616889943   0.17678684090653574   0.4168603844028424   0.7913481699521926   0.5233260639731732   0.6067652342687194   0.470994905056687   0.734465379116517   0.881712120198811   0.34648219008662745   0.5554563816004431   0.8541612884034909   0.4142688249056975   0.7191949652201381   0.45472675614516095   0.10094260357449289   0.218751823365001   0.8702010606631241   0.07359070660535184   0.8001464585233871   0.017254758029190492   0.9046133960897387   0.8869810334680748   0.876723226481039   0.7790455018602911   0.7278265551832028   0.4701206490652324   0.08537505652884635   0.25571943788711793   0.12106132091448349   0.9991257440085454   0.3509096774123293   0.3740073176883069   0.774579130827856   0.44366936240810234   0.4967483890088384   0.9597384927826094   0.05538416560771794   0.9889426062629414   0.3958057854343455   0.7409866694176084   0.18518310494459386   0.9153518996575896   0.5956593269109585   0.723731911388418   0.2805697088548552   0.028370866189514763   0.7189361004299195   0.9446864095281269   0.5527431536716524   0.5582502171242824   0.6335610439010732   0.688966971641009   0.43168183275716887
0.559124473115737   0.2826513664887438   0.314959653952702   0.6571027019293129   0.11545511070763469   0.7859029774799053   0.35522116117009256   0.6017185363215949   0.12651250444469328   0.39009719204555987   0.6142344917524841   0.416535431377001   0.21116060478710375   0.7944378651346015   0.8905025803640663   0.13596572252214575   0.18278973859758899   0.075501764704682   0.9458161708359394   0.5832225688504934   0.6245395214733066   0.44194072080360886   0.25684919919493043   0.15154073609332452   0.06541504835756956   0.1592893543148651   0.9418895452422285   0.4944380341640117   0.9499599376499349   0.3733863768349597   0.5866683840721358   0.8927194978424169   0.8234474332052416   0.9832891847893999   0.9724338923196517   0.47618406646541583   0.6122868284181379   0.18885131965479834   0.08193131195558548   0.3402183439432701   0.42949708982054885   0.11334955495011635   0.1361151411196461   0.7569957750927767   0.8049575683472423   0.6714088341465074   0.8792659419247156   0.6054550389994522   0.7395425199896727   0.5121194798316424   0.9373763966824872   0.11101700483544043   0.7895825823397379   0.13873310299668268   0.3507080126103513   0.21829750699302355   0.9661351491344963   0.15544391820728284   0.37827412029069957   0.7421134405276077   0.3538483207163584   0.9665925985524845   0.29634280833511406   0.4018950965843376
0.9243512308958096   0.8532430436023681   0.160227667215468   0.6448993214915609   0.11939366254856727   0.18183420945586068   0.28096172529075236   0.03944428249210875   0.37985114255889457   0.6697147296242183   0.3435853286082652   0.9284272776566683   0.5902685602191567   0.5309816266275357   0.992877315997914   0.7101297706636448   0.6241334110846605   0.3755377084202528   0.6146031957072143   0.968016330136037   0.270285090368302   0.40894510986776833   0.3182603873721003   0.5661212335516994   0.34593385947249244   0.5557020662654002   0.15803272015663228   0.9212219120601386   0.22654019692392516   0.37386785680953943   0.8770709948658799   0.8817776295680299   0.8466890543650306   0.7041531271853212   0.5334856662576147   0.9533503519113615   0.2564204941458739   0.1731715005577855   0.5406083502597008   0.24322058124771673   0.6322870830612135   0.7976337921375327   0.9260051545524864   0.2752042511116797   0.36200199269291145   0.3886886822697644   0.6077447671803862   0.7090830175599802   0.016068133220419018   0.8329866160043642   0.4497120470237539   0.7878611054998417   0.7895279362964939   0.45911875919482475   0.572641052157874   0.9060834759318118   0.9428388819314633   0.7549656320095036   0.03915538590025925   0.9527331240204504   0.6864183877855894   0.5817941314517181   0.4985470356405584   0.7095125427727337
0.0541313047243759   0.7841603393141855   0.5725418810880719   0.43430829166105395   0.6921293120314644   0.3954716570444211   0.9647971139076857   0.7252252741010737   0.6760611788110454   0.5624850410400569   0.5150850668839319   0.9373641686012321   0.8865332425145516   0.10336628184523211   0.9424440147260579   0.03128069266942027   0.9436943605830883   0.3484006498357285   0.9032886288257986   0.0785475686489699   0.257275972797499   0.7666065183840104   0.4047415931852402   0.36903502587623627   0.20314466807312306   0.9824461790698249   0.8321997120971683   0.9347267342151823   0.5110153560416586   0.5869745220254038   0.8674025981894825   0.20950146011410853   0.8349541772306132   0.024489480985346902   0.3523175313055506   0.2721372915128764   0.9484209347160616   0.9211231991401148   0.4098735165794927   0.24085659884345614   0.004726574132973328   0.5727225493043863   0.506584887753694   0.16230903019448623   0.7474506013354744   0.806116030920376   0.10184329456845385   0.79327400431825   0.5443059332623513   0.8236698518505511   0.2696435824712856   0.8585472701030676   0.03329057722069269   0.23669532982514727   0.40224098428180316   0.6490458099889591   0.1983363999900795   0.21220584883980037   0.04992345297625258   0.37690851847608275   0.24991546527401784   0.2910826496996856   0.6400499363967599   0.1360519196326266
0.24518889114104453   0.7183601003952993   0.1334650486430658   0.9737428894381404   0.49773828980557017   0.9122440694749233   0.03162175407461195   0.1804688851198904   0.9534323565432188   0.08857421762437229   0.7619781716033264   0.3219216150168227   0.9201417793225262   0.851878887799225   0.35973718732152316   0.6728758050278636   0.7218053793324467   0.6396730389594246   0.3098137343452706   0.29596728655178084   0.47188991405842884   0.34859038925973906   0.6697637979485107   0.15991536691915423   0.22670102291738428   0.6302302888644398   0.5362987493054449   0.18617247748101387   0.7289627331118141   0.7179862193895165   0.504676995230833   0.005703592361123463   0.7755303765685954   0.6294120017651441   0.7426988236275066   0.6837819773443008   0.8553885972460692   0.7775331139659191   0.38296163630598345   0.010906172316437177   0.13358321791362252   0.13786007500649447   0.07314790196071287   0.7149388857646564   0.6616933038551936   0.7892696857467554   0.40338410401220215   0.5550235188455022   0.4349922809378094   0.15903939688231566   0.8670853547067573   0.36885104136448826   0.7060295478259953   0.44105317749279926   0.3624083594759243   0.3631474490033648   0.9304991712573999   0.8116411757276552   0.6197095358484177   0.679365471659064   0.07511057401133077   0.03410806176173605   0.23674789954243425   0.6684592993426269
0.9415273560977082   0.8962479867552415   0.16359999758172136   0.9535204135779706   0.27983405224251456   0.10697830100848617   0.7602158935695192   0.3984968947324684   0.8448417713047052   0.9479389041261705   0.893130538862762   0.02964585336798013   0.1388122234787099   0.5068857266333713   0.5307221793868376   0.6664984043646153   0.20831305222130994   0.6952445509057161   0.9110126435384199   0.9871329327055512   0.13320247820997916   0.66113648914398   0.6742647439959857   0.31867363336292437   0.19167512211227092   0.7648885023887385   0.5106647464142643   0.36515321978495385   0.9118410698697563   0.6579102013802522   0.7504488528447452   0.9666563250524854   0.06699929856505121   0.7099712972540818   0.8573183139819832   0.9370104716845054   0.9281870750863414   0.20308557062071053   0.3265961345951456   0.27051206731988997   0.7198740228650314   0.5078410197149944   0.41558349105672565   0.2833791346143387   0.5866715446550522   0.8467045305710144   0.74131874706074   0.9647055012514144   0.39499642254278133   0.08181602818227594   0.23065400064647562   0.5995522814664606   0.48315535267302495   0.42390582680202366   0.4802051478017305   0.6328959564139751   0.41615605410797374   0.7139345295479419   0.6228868338197473   0.6958854847294698   0.4879689790216324   0.5108489589272314   0.2962906992246018   0.4253734174095798
0.768094956156601   0.0030079392122368633   0.8807072081678761   0.14199428279524104   0.18142341150154878   0.15630340864122247   0.13938846110713615   0.17728878154382668   0.7864269889587675   0.07448738045894651   0.9087344604606605   0.5777365000773662   0.3032716362857425   0.6505815536569228   0.42852931265893   0.9448405436633911   0.8871155821777688   0.936647024108981   0.8056424788391827   0.24895505893392134   0.39914660315613637   0.4257980651817497   0.509351779614581   0.8235816415243415   0.6310516469995354   0.4227901259695128   0.6286445714467048   0.6815873587291005   0.44962823549798664   0.2664867173282904   0.4892561103395687   0.5042985771852738   0.6632012465392192   0.19199933686934384   0.5805216498789082   0.9265620771079077   0.35992961025347664   0.541417783212421   0.15199233721997812   0.9817215334445166   0.4728140280757079   0.60477075910344   0.3463498583807954   0.7327664745105953   0.0736674249195715   0.1789726939216903   0.8369980787662145   0.9091848329862537   0.4426157779200361   0.7561825679521774   0.2083535073195096   0.22759747425715318   0.9929875424220495   0.4896958506238871   0.7190973969799409   0.7232988970718793   0.3297862958828303   0.29769651375454326   0.1385757471010328   0.7967368199639716   0.9698566856293537   0.7562787305421222   0.9865834098810546   0.815015286519455
0.4970426575536458   0.15150797143868228   0.6402335515002593   0.08224881200885974   0.4233752326340743   0.972535277516992   0.8032354727340448   0.173063979022606   0.9807594547140381   0.2163527095648145   0.5948819654145352   0.9454665047654528   0.9877719122919887   0.7266568589409274   0.8757845684345942   0.22216760769357347   0.6579856164091583   0.42896034518638415   0.7372088213335615   0.42543078772960186   0.6881289307798046   0.6726816146442619   0.7506254114525068   0.6104155012101469   0.19108627322615887   0.5211736432055796   0.11039185995224754   0.5281666892012871   0.7677110405920846   0.5486383656885876   0.30715638721820276   0.35510271017868106   0.7869515858780464   0.33228565612377314   0.7122744218036676   0.40963620541322826   0.7991796735860578   0.6056287971828457   0.8364898533690733   0.1874685977196548   0.1411940571768994   0.17666845199646158   0.09928103203551195   0.762037809990053   0.45306512639709473   0.5039868373521996   0.34865562058300514   0.15162230877990612   0.2619788531709359   0.98281319414662   0.23826376063075763   0.6234556195786191   0.4942678125788513   0.4341748284580324   0.9311073734125549   0.26835290939993794   0.7073162267008049   0.10188917233425927   0.21883295160888724   0.8587167039867097   0.9081365531147472   0.4962603751514135   0.3823430982398139   0.6712481062670549
0.7669424959378477   0.31959192315495194   0.2830620662043019   0.909210296277002   0.31387736954075296   0.8156050858027523   0.9344064456212967   0.7575879874970959   0.051898516369817106   0.8327918916561322   0.6961426849905391   0.1341323679184768   0.5576307037909658   0.3986170631980998   0.7650353115779843   0.8657794585185389   0.850314477090161   0.29672789086384055   0.546202359969097   0.007062754531829129   0.9421779239754139   0.800467515712427   0.16385926172928314   0.3358146482647742   0.17523542803756614   0.48087559255747503   0.8807971955249813   0.42660435198777225   0.8613580584968131   0.6652705067547228   0.9463907499036844   0.6690163644906764   0.8094595421269961   0.8324786150985906   0.25024806491314533   0.5348839965721995   0.25182883833603026   0.4338615519004907   0.48521275333516106   0.6691045380536608   0.40151436124586926   0.13713366103665012   0.9390103933660641   0.6620417835218316   0.4593364372704554   0.3366661453242231   0.7751511316367808   0.32622713525705743   0.2841010092328892   0.8557905527667481   0.8943539361117997   0.8996227832692851   0.4227429507360761   0.1905200460120253   0.9479631862081153   0.2306064187786088   0.61328340860908   0.35804143091343477   0.6977151212949699   0.6957224222064092   0.3614545702730498   0.9241798790129441   0.2125023679598088   0.026617884152748454
0.9599402090271805   0.7870462179762939   0.2734919745937448   0.36457610063091683   0.5006037717567251   0.45038007265207086   0.4983408429569639   0.03834896537385942   0.21650276252383585   0.5945895198853228   0.6039869068451642   0.13872618210457424   0.7937598117877598   0.4040694738732975   0.6560237206370491   0.9081197633259654   0.18047640317867977   0.04602804295986272   0.9583085993420791   0.21239734111955624   0.81902183290563   0.12184816394691864   0.7458062313822703   0.1857794569668078   0.8590816238784496   0.3348019459706247   0.4723142567885255   0.8212033563358909   0.35847785212172445   0.8844218733185538   0.9739734138315617   0.7828543909620316   0.14197508959788857   0.28983235343323105   0.3699865069863974   0.6441282088574573   0.3482152778101288   0.8857628795599336   0.7139627863493484   0.7360084455314918   0.16773887463144904   0.8397348366000709   0.7556541870072693   0.5236111044119356   0.348717041725819   0.7178866726531522   0.009847955624998956   0.3378316474451278   0.4896354178473695   0.3830847266825275   0.5375336988364734   0.5166282911092368   0.13115756572564508   0.49866285336397365   0.5635602850049118   0.7337739001472053   0.9891824761277564   0.20883049993074262   0.19357377801851441   0.08964569128974798   0.6409671983176277   0.32306762037080905   0.47961099166916604   0.3536372457582561
0.4732283236861786   0.48333278377073824   0.7239568046618968   0.8300261413463206   0.12451128196035961   0.7654461111175861   0.7141088490368979   0.49219449390119274   0.6348758641129901   0.38236138443505857   0.17657515020042439   0.9755662027919559   0.503718298387345   0.8836985310710849   0.6130148651955125   0.2417923026447506   0.5145358222595886   0.6748680311403422   0.41944108717699813   0.15214661135500263   0.8735686239419609   0.3518004107695332   0.9398300955078321   0.7985093655967465   0.4003403002557822   0.868467626998795   0.21587329084593535   0.968483224250426   0.2758290182954226   0.10302151588120892   0.5017644418090376   0.47628873034923325   0.6409531541824325   0.7206601314461504   0.32518929160861315   0.5007225275572773   0.13723485579508746   0.8369616003750655   0.7121744264131006   0.25893022491252676   0.6226990335354989   0.1620935692347232   0.29273333923610245   0.10678361355752411   0.749130409593538   0.81029315846519   0.3529032437282703   0.3082742479607776   0.3487901093377558   0.941825531466395   0.137029952882335   0.33979102371035164   0.07296109104233318   0.8388040155851861   0.6352655110732974   0.8635022933611184   0.4320079368599007   0.11814388413903575   0.31007621946468433   0.362779765803841   0.29477308106481326   0.28118228376397025   0.5979017930515838   0.1038495408913143
0.6720740475293143   0.11908871452924706   0.30516845381548136   0.9970659273337902   0.9229436379357763   0.30879555606405706   0.952265210087211   0.6887916793730126   0.5741535285980205   0.36697002459766204   0.815235257204876   0.349000655662661   0.5011924375556873   0.5281660090124759   0.17996974613157854   0.48549836230154253   0.06918450069578663   0.41002212487344014   0.8698935266668942   0.1227185964977015   0.7744114196309734   0.1288398411094699   0.2719917336153104   0.018869055606387193   0.10233737210165907   0.009751126580222834   0.9668232797998291   0.02180312827259699   0.17939373416588275   0.7009555705161657   0.01455806971261805   0.3330114488995844   0.6052402055678623   0.33398554591850377   0.19932281250774203   0.9840107932369234   0.10404776801217493   0.8058195369060278   0.019353066376163477   0.4985124309353809   0.0348632673163883   0.3957974120325877   0.14945953970926928   0.3757938344376794   0.2604518476854149   0.26695757092311784   0.8774678060939589   0.3569247788312922   0.15811447558375585   0.25720644434289497   0.9106445262941298   0.3351216505586952   0.9787207414178731   0.5562508738267292   0.8960864565815118   0.002110201659110814   0.37348053585001084   0.22226532790822545   0.6967636440737697   0.018099408422187362   0.26943276783783593   0.4164457910021976   0.6774105776976063   0.5195869774868065
0.23456950052144762   0.020648378969609867   0.527951037988337   0.14379314304912708   0.9741176528360327   0.753690808046492   0.6504832318943781   0.7868683642178349   0.8160031772522769   0.49648436370359705   0.7398387056002483   0.45174671365913965   0.8372824358344038   0.9402334898768678   0.8437522490187366   0.4496365120000288   0.4638018999843929   0.7179681619686424   0.14698860494496682   0.4315371035778415   0.19436913214655702   0.30152237096644485   0.4695780272473606   0.911950126091035   0.9597996316251094   0.280873991996835   0.9416269892590237   0.7681569830419079   0.9856819787890767   0.5271831839503429   0.29114375736464554   0.981288618824073   0.16967880153679984   0.03069882024674587   0.5513050517643973   0.5295419051649335   0.3323963657023961   0.09046533036987803   0.7075528027456607   0.07990539316490462   0.8685944657180031   0.3724971684012356   0.5605641978006939   0.6483682895870632   0.6742253335714461   0.07097479743479078   0.09098617055333327   0.7364181634960282   0.7144257019463367   0.7901008054379558   0.14935918129430967   0.9682611804541202   0.72874372315726   0.2629176214876129   0.8582154239296641   0.9869725616300471   0.5590649216204602   0.23221880124086702   0.3069103721652669   0.45743065646511366   0.22666855591806404   0.141753470870989   0.5993575694196063   0.3775252633002091
0.35807409020006087   0.7692563024697534   0.03879337161891237   0.7291569737131459   0.6838487566286148   0.6982815050349626   0.9478072010655791   0.9927388102171177   0.9694230546822781   0.9081806995970068   0.7984480197712694   0.024477629762997555   0.24067933152501808   0.6452630781093939   0.9402325958416053   0.03750506813295043   0.681614409904558   0.41304427686852685   0.6333222236763384   0.5800744116678368   0.45494585398649395   0.27129080599753785   0.033964654256732174   0.20254914836762766   0.09687176378643304   0.5020345035277844   0.9951712826378198   0.47339217465448175   0.41302300715781826   0.8037529984928219   0.0473640815722407   0.480653364437364   0.4435999524755402   0.8955722988958151   0.24891606180097126   0.45617573467436645   0.2029206209505221   0.2503092207864212   0.30868346595936597   0.418670666541416   0.5213062110459642   0.8372649439178943   0.6753612422830275   0.8385962548735792   0.06636035705947022   0.5659741379203564   0.6413965880262954   0.6360471065059516   0.9694885932730372   0.06393963439257197   0.6462253053884756   0.16265493185146984   0.5564655861152189   0.2601866358997501   0.5988612238162349   0.6820015674141059   0.1128656336396787   0.36461433700393503   0.3499451620152636   0.22582583273973938   0.9099450126891566   0.11430511621751382   0.04126169605589766   0.8071551661983234
0.3886388016431924   0.2770401722996195   0.3659004537728701   0.9685589113247441   0.32227844458372223   0.7110660343792631   0.7245038657465747   0.33251180481879256   0.352789851310685   0.6471263999866911   0.07827856035809912   0.16985687296732271   0.7963242651954662   0.386939764086941   0.47941733654186425   0.4878553055532169   0.6834586315557875   0.022325427083005955   0.1294721745266006   0.2620294728134775   0.7735136188666308   0.9080203108654922   0.08821047847070294   0.4548743066151541   0.3848748172234384   0.6309801385658727   0.7223100246978328   0.48631539529040996   0.06259637263971618   0.9199141041866096   0.9978061589512581   0.15380359047161743   0.7098065213290311   0.2727877041999185   0.919527598593159   0.9839467175042947   0.913482256133565   0.8858479401129775   0.4401102620512948   0.49609141195107787   0.23002362457777756   0.8635225130299715   0.3106380875246942   0.2340619391376004   0.4565100057111467   0.9555022021644795   0.22242760905399125   0.7791876325224463   0.0716351884877083   0.3245220635986068   0.5001175843561584   0.29287223723203637   0.009038815847992127   0.40460795941199723   0.5023114254049003   0.13906864676041894   0.299232294518961   0.13182025521207874   0.5827838268117412   0.1551219292561242   0.385750038385396   0.24597231509910122   0.14267356476044646   0.6590305173050464
0.15572641380761845   0.38244980206912965   0.8320354772357523   0.42496857816744593   0.6992164080964718   0.4269475999046502   0.609607868181761   0.6457809456449997   0.6275812196087635   0.1024255363060434   0.10949028382560262   0.3529087084129633   0.6185424037607713   0.6978175768940461   0.6071788584207023   0.21384006165254435   0.3193101092418103   0.5659973216819674   0.02439503160896108   0.05871813239642013   0.9335600708564143   0.3200250065828662   0.8817214668485146   0.3996876150913738   0.7778336570487958   0.9375752045137365   0.04968598961276233   0.9747190369239278   0.07861724895232411   0.5106276046090863   0.4400781214310013   0.3289380912789282   0.4510360293435607   0.40820206830304295   0.33058783760539867   0.9760293828659649   0.8324936255827894   0.7103844914089967   0.7234089791846964   0.7621893212134205   0.513183516340979   0.14438716972702936   0.6990139475757352   0.7034711888170004   0.5796234454845647   0.8243621631441631   0.8172924807272206   0.30378357372562664   0.8017897884357689   0.8867869586304266   0.7676064911144583   0.32906453680169884   0.7231725394834447   0.37615935402134026   0.327528369683457   0.00012644552277063298   0.2721365101398841   0.9679572857182973   0.9969405320780583   0.02409706265680572   0.4396428845570947   0.2575727943093006   0.273531552893362   0.26190774144338513
0.9264593682161157   0.11318562458227122   0.5745176053176267   0.5584365526263847   0.34683592273155095   0.28882346143810805   0.7572251245904061   0.25465297890075805   0.5450461342957821   0.40203650280768144   0.9896186334759478   0.9255884420990592   0.8218735948123373   0.025877148786341182   0.6620902637924907   0.9254619965762886   0.5497370846724533   0.05791986306804384   0.6651497317144324   0.9013649339194829   0.11009420011535856   0.8003470687587433   0.3916181788210704   0.6394571924760978   0.18363483189924287   0.6871614441764721   0.8171005735034437   0.08102063984971301   0.836798909167692   0.398337982738364   0.05987544891303759   0.826367660948955   0.2917527748719098   0.9963014799306825   0.07025681543708982   0.9007792188498958   0.4698791800595724   0.9704243311443413   0.4081665516445991   0.9753172222736071   0.9201420953871191   0.9125044680762975   0.7430168199301667   0.07395228835412421   0.8100478952717606   0.11215739931755425   0.35139864110909624   0.4344950958780265   0.6264130633725177   0.4249959551410822   0.5342980676056526   0.35347445602831346   0.7896141542048258   0.026657972402718177   0.474422618692615   0.5271067950793585   0.497861379332916   0.030356492472035618   0.4041658032555252   0.6263275762294628   0.02798219927334358   0.059932161327694244   0.9959992516109261   0.6510103539558557
0.10784010388622443   0.1474276932513967   0.25298243168075946   0.5770580656017315   0.29779220861446387   0.035270293933842456   0.9015837905716632   0.14256296972370502   0.6713791452419462   0.6102743387927603   0.3672857229660106   0.7890885136953916   0.8817649910371204   0.5836163663900421   0.8928631042733957   0.2619817186160331   0.38390361170420434   0.5532598739180065   0.48869730101787046   0.6356541423865703   0.3559214124308608   0.4933277125903122   0.49269804940694434   0.9846437884307145   0.24808130854463634   0.3459000193389155   0.23971561772618488   0.4075857228289831   0.9502890999301725   0.31062972540507305   0.33813182715452167   0.26502275310527806   0.2789099546882263   0.7003553866123128   0.970846104188511   0.4759342394098865   0.39714496365110596   0.1167390202222707   0.07798299991511547   0.2139525207938534   0.01324135194690158   0.5634791463042642   0.589285698897245   0.5782983784072832   0.6573199395160408   0.07015143371395198   0.09658764949030069   0.5936545899765685   0.40923863097140445   0.7242514143750365   0.8568720317641157   0.18606886714758544   0.458949531041232   0.4136216889699634   0.5187402046095941   0.9210461140423074   0.18003957635300566   0.7132663023576505   0.547894100421083   0.4451118746324209   0.7828946127018998   0.5965272821353799   0.46991110050596757   0.2311593538385675
0.7696532607549982   0.03304813583111568   0.8806254016087225   0.6528609754312844   0.11233332123895733   0.9628967021171637   0.7840377521184219   0.05920638545471587   0.7030946902675529   0.23864528774212726   0.927165720354306   0.8731375183071304   0.2441451592263209   0.8250235987721639   0.4084255157447119   0.9520914042648231   0.06410558287331526   0.11175729641451328   0.8605314153236289   0.5069795296324021   0.28121097017141555   0.5152300142791334   0.39062031481766135   0.27582017579383467   0.5115577094164174   0.4821818784480177   0.5099949132089387   0.6229592003625503   0.3992243881774601   0.519285176330854   0.725957161090517   0.5637528149078344   0.6961296979099072   0.28063988858872674   0.7987914407362109   0.690615296600704   0.4519845386835863   0.4556162898165629   0.39036592499149897   0.7385238923358809   0.38787895581027104   0.3438589934020496   0.52983450966787   0.23154436270347875   0.10666798563885548   0.8286289791229162   0.1392141948502087   0.9557241869096441   0.5951102762224381   0.34644710067489853   0.6292192816412698   0.33276498654709386   0.19588588804497795   0.8271619243440446   0.903262120550753   0.7690121716392595   0.4997561901350707   0.5465220357553178   0.10447067981454204   0.0783968750385555   0.047771651451484425   0.0909057459387549   0.7141047548230431   0.3398729827026746
0.6598926956412134   0.7470467525367053   0.18427024515517307   0.10832861999919584   0.553224710002358   0.918417773413789   0.04505605030496438   0.15260443308955174   0.9581144337799199   0.5719706727388906   0.4158367686636945   0.8198394465424579   0.7622285457349419   0.744808748394846   0.5125746481129415   0.05082727490319842   0.26247235559987125   0.19828671263952824   0.4081039682983995   0.972430399864643   0.2147007041483868   0.10738096670077334   0.6939992134753564   0.6325574171619683   0.5548080085071734   0.360334214164068   0.5097289683201833   0.5242287971627725   0.001583298504815482   0.44191644075027897   0.464672918015219   0.37162436407322075   0.04346886472489559   0.8699457680113885   0.048836149351524465   0.5517849175307629   0.28124031898995366   0.1251370196165424   0.5362615012385828   0.5009576426275645   0.018767963390082413   0.9268503069770141   0.1281575329401834   0.5285272427629215   0.8040672592416956   0.8194693402762409   0.43415831946482697   0.8959698256009532   0.2492592507345222   0.4591351261121728   0.9244293511446436   0.37174102843818074   0.24767595222970673   0.01721868536189379   0.45975643312942466   0.00011666436495997266   0.20420708750481112   0.14727291735050538   0.4109202837779002   0.4483317468341971   0.9229667685148575   0.022135897733962982   0.8746587825393173   0.9473741042066326
0.904198805124775   0.09528559075694884   0.7465012495991339   0.4188468614437111   0.10013154588307946   0.275816250480708   0.3123429301343069   0.5228770358427578   0.8508722951485572   0.8166811243685352   0.38791357898966333   0.1511360074045771   0.6031963429188505   0.7994624390066415   0.9281571458602387   0.15101934303961712   0.3989892554140394   0.6521895216561361   0.5172368620823384   0.70268759620542   0.4760224868991819   0.6300536239221731   0.6425780795430212   0.7553134919987874   0.5718236817744069   0.5347680331652243   0.8960768299438873   0.33646663055507636   0.4716921358913274   0.25895178268451624   0.5837338998095803   0.8135895947123185   0.6208198407427702   0.442270658315981   0.19582032081991702   0.6624535873077414   0.0176234978239196   0.6428082193093395   0.26766317495967834   0.5114342442681243   0.6186342424098802   0.9906186976532034   0.7504263128773399   0.8087466480627042   0.14261175551069827   0.36056507373103025   0.10784823333431873   0.05343315606391684   0.5707880737362914   0.8257970405658059   0.21177140339043146   0.7169665255088404   0.099095937844964   0.5668452578812897   0.6280375035808511   0.9033769307965219   0.4782760971021939   0.12457459956530875   0.4322171827609341   0.24092334348878053   0.46065259927827423   0.48176638025596924   0.16455400780125576   0.7294890992206562
0.8420183568683941   0.49114768260276587   0.4141276949239159   0.920742451157952   0.6994066013576958   0.1305826088717356   0.3062794615895971   0.8673092950940351   0.1286185276214044   0.30478556830592957   0.09450805819916568   0.15034276958519463   0.02952258977644042   0.7379403104246398   0.46647055461831455   0.2469658387886727   0.5512464926742465   0.6133657108593311   0.03425337185738042   0.0060424952998921685   0.09059389339597232   0.13159933060336185   0.8696993640561247   0.27655339607923596   0.24857553652757824   0.640451648000596   0.4555716691322088   0.355810944921284   0.5491689351698824   0.5098690391288604   0.1492922075426117   0.48850164982724886   0.42055040754847806   0.20508347082293082   0.054784149343446005   0.33815888024205426   0.3910278177720376   0.46714316039829096   0.5883135947251315   0.09119304145338154   0.839781325097791   0.8537774495389598   0.554060222867751   0.08515054615348938   0.7491874317018187   0.722178118935598   0.6843608588116263   0.8085971500742535   0.5006118951742404   0.08172647093500207   0.22878918967941758   0.4527862051529694   0.951442960004358   0.5718574318061417   0.0794969821368059   0.9642845553257205   0.53089255245588   0.36677396098321086   0.024712832793359892   0.6261256750836663   0.13986473468384236   0.8996308005849198   0.43639923806822845   0.5349326336302848
0.30008340958605134   0.04585335104595999   0.8823390152004774   0.4497820874767954   0.5508959778842326   0.3236752321103619   0.197978156388851   0.641184937402542   0.050284082709992135   0.24194876117535988   0.9691889667094334   0.18839873224957254   0.09884112270563412   0.6700913293692182   0.8896919845726275   0.22411417692385197   0.5679485702497541   0.30331736838600737   0.8649791517792677   0.5979885018401857   0.4280838355659118   0.4036865678010875   0.4285799137110392   0.06305586820990088   0.12800042597986044   0.3578332167551275   0.5462408985105618   0.6132737807331055   0.5771044480956279   0.03415798464476556   0.3482627421217108   0.9720888433305636   0.5268203653856357   0.7922092234694057   0.37907377541227744   0.783690111080991   0.4279792426800016   0.12211789410018746   0.4893817908396499   0.559575934157139   0.8600306724302474   0.81880052571418   0.6244026390603823   0.9615874323169533   0.4319468368643357   0.4151139579130926   0.19582272534934306   0.8985315641070525   0.3039464108844752   0.05728074115796507   0.6495818268387812   0.285257783373947   0.7268419627888474   0.02312275651319951   0.30131908471707036   0.31316894004338347   0.20002159740321165   0.23091353304379383   0.922245309304793   0.5294788289623925   0.77204235472321   0.10879563894360637   0.43286351846514304   0.9699028948052535
0.9120116822929626   0.2899951132294263   0.8084608794047607   0.00831546248830009   0.4800648454286269   0.8748811553163337   0.6126381540554178   0.10978389838124761   0.17611843454415166   0.8176004141583687   0.9630563272166365   0.8245261150073006   0.4492764717553043   0.7944776576451692   0.6617372424995661   0.5113571749639171   0.24925487435209262   0.5635641246013753   0.7394919331947731   0.9818783460015247   0.47721251962888256   0.45476848565776895   0.3066284147296301   0.011975451196271178   0.56520083733592   0.16477337242834264   0.4981675353248693   0.0036599887079710866   0.0851359919072931   0.2898922171120089   0.8855293812694516   0.8938760903267234   0.9090175573631414   0.47229180295364026   0.9224730540528151   0.06934997531942289   0.45974108560783716   0.6778141453084711   0.26073581155324893   0.5579928003555058   0.21048621125574452   0.1142500207070958   0.5212438783584757   0.5761144543539811   0.733273691626862   0.6594815350493268   0.21461546362884568   0.5641390031577099   0.16807285429094196   0.4947081626209842   0.7164479283039763   0.5604790144497389   0.08293686238364885   0.2048159455089753   0.8309185470345247   0.6666029241230154   0.17391930502050743   0.732524142555335   0.9084454929817097   0.5972529488035925   0.7141782194126702   0.05470999724686392   0.6477096814284607   0.03926014844808673
0.5036920081569257   0.9404599765397681   0.12646580306998498   0.4631456940941056   0.7704183165300638   0.28097844149044127   0.9118503394411394   0.8990066909363956   0.6023454622391219   0.786270278869457   0.19540241113716295   0.3385276764866568   0.5194085998554729   0.5814543333604817   0.36448386410263817   0.6719247523636415   0.3454892948349656   0.8489301908051468   0.4560383711209285   0.07467180356004895   0.6313110754222954   0.7942201935582828   0.8083286896924677   0.03541165511196222   0.12761906726536956   0.8537602170185147   0.6818628866224827   0.5722659610178567   0.35720075073530577   0.5727817755280734   0.7700125471813435   0.6732592700814609   0.7548552884961839   0.7865114966586163   0.5746101360441805   0.33473159359480414   0.23544668864071094   0.20505716329813461   0.2101262719415423   0.6628068412311627   0.8899573938057453   0.3561269724929879   0.7540879008206138   0.5881350376711137   0.25864631838345004   0.5619067789347051   0.9457592111281461   0.5527233825591515   0.13102725111808047   0.7081465619161905   0.2638963245056633   0.9804574215412949   0.7738265003827747   0.13536478638811708   0.4938837773243199   0.307198151459834   0.018971211886590775   0.3488532897295007   0.9192736412801393   0.9724665578650298   0.7835245232458798   0.1437961264313661   0.709147369338597   0.30965971663386715
0.8935671294401345   0.7876691539383782   0.9550594685179833   0.7215246789627534   0.6349208110566844   0.22576237500367305   0.009300257389837172   0.16880129640360184   0.503893559938604   0.5176158130874826   0.7454039328841738   0.18834387486230691   0.7300670595558293   0.3822510266993655   0.251520155559854   0.881145723402473   0.7110958476692385   0.033397736969864804   0.33224651427971463   0.9086791655374431   0.9275713244233587   0.8896016105384987   0.6230991449411176   0.599019448903576   0.03400419498322416   0.10193245660012053   0.6680396764231343   0.8774947699408226   0.3990833839265397   0.8761700815964475   0.6587394190332971   0.7086934735372208   0.8951898239879358   0.3585542685089649   0.9133354861491233   0.5203495986749138   0.16512276443210647   0.9763032418095994   0.6618153305892693   0.6392038752724409   0.454026916762868   0.9429055048397346   0.32956881630955465   0.7305247097349978   0.5264555923395093   0.05330389430123586   0.7064696713684371   0.13150526083142183   0.4924513973562852   0.9513714377011153   0.038429994945302755   0.25401049089059924   0.09336801342974545   0.07520135610466787   0.3796905759120056   0.5453170173533785   0.1981781894418097   0.716647087595703   0.4663550897628823   0.024967418678464626   0.03305542500970324   0.7403438457861036   0.804539759173613   0.3857635434060237
0.5790285082468353   0.797438340946369   0.47497094286405833   0.6552388336710259   0.05257291590732594   0.7441344466451332   0.7685012714956212   0.5237335728396041   0.5601215185510408   0.7927630089440179   0.7300712765503184   0.2697230819490048   0.4667535051212953   0.71756165283935   0.3503807006383129   0.7244060645956264   0.2685753156794856   0.0009145652436469969   0.8840256108754306   0.6994386459171618   0.2355198906697824   0.2605707194575434   0.07948585170181759   0.313675102511138   0.6564913824229471   0.46313237851117434   0.6045149088377593   0.6584362688401121   0.6039184665156212   0.7189979318660411   0.836013637342138   0.13470269600050805   0.043796947964580404   0.9262349229220233   0.10594236079181953   0.8649796140515033   0.5770434428432851   0.20867327008267333   0.7555616601535067   0.14057354945587688   0.30846812716379945   0.20775870483902634   0.871536049278076   0.44113490353871515   0.07294823649401705   0.947187985381483   0.7920501975762585   0.12745980102757715   0.4164568540710699   0.48405560687030863   0.1875352887384992   0.46902353218746506   0.8125383875554487   0.7650576750042675   0.35152165139636116   0.334320836186957   0.7687414395908683   0.8388227520822441   0.24557929060454164   0.46934122213545376   0.19169799674758325   0.6301494819995709   0.490017630451035   0.3287676726795769
0.8832298695837838   0.4223907771605445   0.618481581172959   0.8876327691408618   0.8102816330897668   0.47520279177906155   0.8264313835967005   0.7601729681132846   0.39382477901869684   0.991147184908753   0.6388960948582013   0.29114943592581954   0.5812863914632481   0.2260895099044855   0.28737444346184016   0.9568285997388625   0.8125449518723799   0.38726675782224135   0.04179515285729851   0.48748737760340877   0.6208469551247966   0.7571172758226705   0.5517775224062635   0.15871970492383183   0.7376170855410128   0.334726498662126   0.9332959412333045   0.2710869357829701   0.927335452451246   0.8595237068830645   0.10686455763660398   0.5109139676696856   0.5335106734325491   0.8683765219743115   0.46796846277840265   0.21976453174386595   0.952224281969301   0.642287012069826   0.18059401931656247   0.2629359320050034   0.13967933009692124   0.2550202542475846   0.13879886645926395   0.7754485544015947   0.5188323749721246   0.4979029784249141   0.5870213440530004   0.6167288494777629   0.781215289431112   0.1631764797627881   0.6537254028196959   0.34564191369479275   0.8538798369798659   0.30365277287972364   0.546860845183092   0.8347279460251072   0.32036916354731676   0.43527625090541217   0.07889238240468935   0.6149634142812413   0.3681448815780157   0.7929892388355861   0.8982983630881269   0.35202748227623787
0.22846555148109451   0.5379689845880015   0.759499496628863   0.5765789278746432   0.7096331765089698   0.04006600616308739   0.1724781525758625   0.9598500783968803   0.9284178870778579   0.8768895264002993   0.5187527497561666   0.6142081647020875   0.074538050097992   0.5732367535205757   0.9718919045730746   0.7794802186769803   0.7541688865506753   0.13796050261516352   0.8929995221683852   0.16451680439573896   0.3860240049726595   0.3449712637795774   0.9947011590802584   0.8124893221195011   0.157558453491565   0.8070022791915759   0.2352016624513954   0.23591039424485793   0.44792527698259516   0.7669362730284884   0.06272350987553288   0.27606031584797763   0.5195073899047372   0.8900467466281892   0.5439707601193663   0.6618521511458901   0.44496933980674525   0.3168099931076135   0.5720788555462918   0.8823719324689099   0.69080045325607   0.17884949049245   0.6790793333779065   0.7178551280731709   0.3047764482834105   0.8338782267128726   0.6843781742976481   0.9053658059536698   0.14721799479184552   0.0268759475212968   0.4491765118462528   0.6694554117088118   0.6992927178092504   0.25993967449280836   0.3864530019707199   0.39339509586083427   0.17978532790451313   0.3698929278646192   0.8424822418513536   0.7315429447149442   0.7348159880977679   0.05308293475700571   0.27040338630506183   0.8491710122460343
0.04401553484169788   0.8742334442645557   0.5913240529271553   0.1313158841728634   0.7392390865582874   0.04035521755168307   0.9069458786295072   0.22595007821919358   0.5920210917664418   0.013479270030386273   0.4577693667832544   0.5564946665103817   0.8927283739571914   0.7535395955375779   0.0713163648125345   0.16309957064954744   0.7129430460526783   0.3836466676729587   0.22883412296118094   0.4315566259346033   0.9781270579549104   0.330563732915953   0.9584307366561191   0.582385613688569   0.9341115231132125   0.4563302886513973   0.36710668372896377   0.45106972951570556   0.19487243655492517   0.4159750710997142   0.4601608050994566   0.22511965129651199   0.6028513447884833   0.4024958010693279   0.0023914383162021956   0.6686249847861303   0.7101229708312919   0.64895620553175   0.9310750735036677   0.5055254141365828   0.9971799247786136   0.2653095378587913   0.7022409505424867   0.07396878820197955   0.019052866823703173   0.9347458049428383   0.7438102138863676   0.49158317451341055   0.08494134371049064   0.478415516291441   0.3767035301574039   0.04051344499770497   0.8900689071555654   0.06244044519172685   0.9165427250579473   0.815393793701193   0.2872175623670821   0.659944644122399   0.9141512867417451   0.1467688089150627   0.5770945915357902   0.010988438590648908   0.9830762132380774   0.6412433947784798
0.5799146667571766   0.7456789007318576   0.2808352626955906   0.5672746065765003   0.5608617999334734   0.8109330957890193   0.537025048809223   0.07569143206308974   0.4759204562229828   0.33251757949757826   0.16032151865181915   0.035177987065384775   0.5858515490674173   0.2700771343058514   0.24377879359387186   0.2197841933641918   0.29863398670033525   0.6101324901834525   0.32962750685212683   0.07301538444912913   0.721539395164545   0.5991440515928036   0.3465512936140494   0.4317719896706493   0.14162472840736837   0.853465150860946   0.06571603091845878   0.864497383094149   0.5807629284738949   0.042532055071926686   0.5286909821092358   0.7888059510310592   0.1048424722509121   0.7100144755743485   0.3683694634574166   0.7536279639656744   0.5189909231834947   0.43993734126849704   0.12459066986354476   0.5338437706014827   0.22035693648315952   0.8298048510850445   0.794963163011418   0.46082838615235355   0.4988175413186145   0.230660799492241   0.44841186939736855   0.029056396481704265   0.35719281291124616   0.377195648631295   0.38269583847890976   0.16455901338755527   0.7764298844373512   0.33466359355936837   0.854004856369674   0.375753062356496   0.6715874121864391   0.6246491179850199   0.4856353929122574   0.6221250983908215   0.15259648900294437   0.18471177671652286   0.3610447230487126   0.08828132778933889
0.9322395525197849   0.3549069256314783   0.5660815600372946   0.6274529416369854   0.4334220112011703   0.12424612613923729   0.1176696906399261   0.5983965451552811   0.07622919828992418   0.7470504775079423   0.7349738521610163   0.43383753176772577   0.29979931385257297   0.4123868839485739   0.8809689957913424   0.058084469411229765   0.6282119016661338   0.787737765963554   0.395333602879085   0.4359593710204082   0.4756154126631895   0.6030259892470312   0.03428887983037238   0.3476780432310693   0.5433758601434047   0.2481190636155529   0.4682073197930777   0.7202251015940839   0.10995384894223435   0.1238729374763156   0.3505376291531516   0.1218285564388029   0.033724650652310166   0.3768224599683733   0.6155637769921353   0.6879910246710771   0.7339253367997371   0.9644355760197995   0.7345947812007929   0.6299065552598473   0.10571343513360335   0.1766978100562454   0.339261178321708   0.19394718423943913   0.6300980224704138   0.5736718208092142   0.3049722984913356   0.8462691410083698   0.08672216232700919   0.3255527571936614   0.8367649786982578   0.12604403941428585   0.9767683133847749   0.20167981971734578   0.4862273495451062   0.0042154829754829475   0.9430436627324646   0.8248573597489725   0.8706635725529709   0.3162244583044059   0.20911832593272747   0.860421783729173   0.13606879135217795   0.6863179030445585
0.10340489079912413   0.6837239736729276   0.79680761303047   0.4923707188051194   0.4733068683287103   0.11005215286371334   0.49183531453913437   0.6461015777967496   0.3865847060017011   0.784499395670052   0.6550703358408765   0.5200575383824637   0.40981639261692626   0.5828195759527062   0.16884298629577027   0.5158420554069808   0.46677272988446156   0.7579622162037338   0.2981794137427993   0.19961759710257493   0.2576544039517341   0.8975404324745608   0.16211062239062138   0.5132996940580165   0.15424951315260998   0.2138164588016332   0.3653030093601514   0.020928975252897032   0.6809426448238998   0.10376430593791987   0.873467694821017   0.37482739745614746   0.29435793882219863   0.3192649102678679   0.21839735898014057   0.8547698590736837   0.8845415462052724   0.7364453343151617   0.049554372684370296   0.33892780366670294   0.4177688163208108   0.978483118111428   0.7513749589415709   0.13931020656412804   0.1601144123690767   0.08094268563686713   0.5892643365509496   0.6260105125061116   0.005864899216466696   0.8671262268352339   0.22396132719079814   0.6050815372532146   0.324922254392567   0.763361920897314   0.3504936323697811   0.23025413979706713   0.030564315570368344   0.4440970106294462   0.1320962733896405   0.3754842807233834   0.14602276936509595   0.7076516763142845   0.08254190070527022   0.03655647705668043
0.7282539530442852   0.7291685582028565   0.33116694176369926   0.8972462704925523   0.5681395406752084   0.6482258725659894   0.7419026052127498   0.2712357579864408   0.5622746414587417   0.7810996457307555   0.5179412780219516   0.6661542207332262   0.2373523870661748   0.01773772483344144   0.1674476456521705   0.43590008093615906   0.20678807149580647   0.5736407142039953   0.03535137226252997   0.06041580021277567   0.0607653021307105   0.8659890378897108   0.9528094715572597   0.02385932315609525   0.3325113490864253   0.1368204796868542   0.6216425297935605   0.12661305266354286   0.7643718084112169   0.4885946071208648   0.8797399245808107   0.8553772946771021   0.2020971669524751   0.7074949613901093   0.36179864655885924   0.1892230739438759   0.9647447798863003   0.6897572365566678   0.19435100090668875   0.7533229930077169   0.7579567083904938   0.11611652235267256   0.15899962864415876   0.6929071927949412   0.6971914062597834   0.2501274844629618   0.20619015708689903   0.6690478696388459   0.364680057173358   0.11330700477610756   0.5845476272933385   0.542434816975303   0.6003082487621412   0.6247123976552428   0.7048077027125278   0.6870575222982009   0.398211081809666   0.9172174362651335   0.3430090561536685   0.49783444835432505   0.43346630192336577   0.2274601997084657   0.14865805524697978   0.7445114553466082
0.6755095935328719   0.11134367735579316   0.989658426602821   0.05160426255166707   0.9783181872730886   0.8612161928928314   0.783468269515922   0.3825563929128212   0.6136381300997306   0.7479091881167238   0.19892064222258346   0.8401215759375181   0.013329881337589458   0.12319679046148105   0.49411293951005575   0.1530640536393171   0.6151187995279234   0.2059793541963475   0.15110388335638722   0.6552296052849921   0.18165249760455765   0.9785191544878817   0.0024458281094074264   0.9107181499383838   0.5061429040716857   0.8671754771320886   0.012787401506586417   0.8591138873867168   0.5278247167985971   0.005959284239257224   0.22931913199066442   0.47655749447389556   0.9141865866988665   0.2580500961225334   0.030398489768080957   0.6364359185363775   0.900856705361277   0.13485330566105236   0.5362855502580253   0.48337186489706035   0.2857379058333537   0.9288739514647049   0.385181666901638   0.8281422596120683   0.10408540822879603   0.950354796976823   0.3827358387922306   0.9174241096736845   0.5979425041571103   0.08317931984473442   0.3699484372856442   0.0583102222869678   0.07011778735851315   0.0772200356054772   0.14062930529497977   0.5817527278130722   0.15593120065964658   0.8191699394829438   0.1102308155268988   0.9453168092766947   0.2550744952983695   0.6843166338218915   0.5739452652688736   0.46194494437963435
0.9693365894650158   0.7554426823571866   0.18876359836723555   0.633802684767566   0.8652511812362198   0.8050878853803636   0.8060277595750049   0.7163785750938815   0.2673086770791095   0.7219085655356291   0.43607932228936075   0.6580683528069137   0.19719088972059634   0.6446885299301519   0.295450016994381   0.07631562499384145   0.04125968906094976   0.8255185904472081   0.1852192014674822   0.13099881571714672   0.7861851937625802   0.14120195662531665   0.6112739361986086   0.6690538713375124   0.8168486042975645   0.38575927426813   0.4225103378313731   0.0352511865699464   0.9515974230613446   0.5806713888877665   0.6164825782563681   0.31887261147606494   0.6842887459822352   0.8587628233521373   0.1804032559670074   0.6608042586691513   0.4870978562616388   0.21407429342198533   0.8849532389726263   0.5844886336753098   0.4458381672006891   0.3885557029747772   0.6997340375051442   0.4534898179581631   0.6596529734381088   0.24735374634946056   0.08846010130653557   0.7844359466206507   0.8428043691405444   0.8615944720813306   0.6659497634751625   0.7491847600507043   0.8912069460791997   0.28092308319356407   0.04946718521879435   0.4303121485746394   0.2069182000969645   0.4221602598414268   0.869063929251787   0.7695078899054881   0.7198203438353257   0.20808596641944144   0.9841106902791605   0.18501925623017826
0.2739821766346366   0.8195302634446643   0.28437665277401636   0.7315294382720151   0.6143292031965278   0.5721765170952037   0.19591655146748077   0.9470934916513645   0.7715248340559835   0.7105820450138731   0.5299667879923182   0.19790873160066014   0.8803178879767838   0.4296589618203091   0.48049960277352394   0.7675965830260207   0.6733996878798193   0.007498701978882286   0.611435673521737   0.9980886931205327   0.9535793440444936   0.7994127355594408   0.6273249832425765   0.8130694368903544   0.6795971674098571   0.9798824721147766   0.3429483304685601   0.08153999861833926   0.06526796421332925   0.4077059550195729   0.1470317790010793   0.1344465069669748   0.29374313015734577   0.6971239100056997   0.617064991008761   0.9365377753663147   0.413425242180562   0.2674649481853907   0.1365653882352371   0.16894119234029387   0.7400255543007427   0.2599662462065084   0.5251297147135001   0.1708524992197612   0.7864462102562491   0.46055351064706757   0.8978047314709237   0.35778306232940676   0.10684904284639198   0.48067103853229093   0.5548564010023637   0.27624306371106755   0.04158107863306273   0.07296508351271803   0.40782462200128433   0.14179655674409272   0.7478379484757169   0.3758411735070183   0.7907596309925233   0.2052587813777781   0.33441270629515496   0.10837622532162762   0.6541942427572862   0.0363175890374842
0.5943871519944123   0.8484099791151193   0.12906452804378607   0.865465089817723   0.8079409417381632   0.3878564684680517   0.23125979657286236   0.5076820274883163   0.7010918988917713   0.9071854299357608   0.6764033955704988   0.2314389637772487   0.6595108202587086   0.8342203464230427   0.26857877356921445   0.08964240703315599   0.9116728717829916   0.4583791729160244   0.47781914257669117   0.8843836256553779   0.5772601654878367   0.35000294759439676   0.823624899819405   0.8480660366178937   0.9828730134934244   0.5015929684792776   0.6945603717756189   0.9826009468001707   0.17493207175526115   0.11373650001122584   0.4633005752027565   0.4749189193118545   0.4738401728634899   0.20655107007546508   0.7868971796322578   0.24347995553460575   0.8143293526047813   0.37233072365242237   0.5183184060630434   0.15383754850144976   0.9026564808217898   0.913951550736398   0.04049926348635222   0.2694539228460719   0.3253963153339532   0.5639486031420011   0.21687436366694726   0.4213878862281782   0.34252330184052876   0.06235563466272363   0.5223139918913283   0.43878693942800745   0.16759123008526763   0.9486191346514978   0.05901341668857179   0.963868020116153   0.6937510572217778   0.7420680645760327   0.272116237056314   0.7203880645815472   0.8794217046169963   0.3697373409236103   0.7537978309932706   0.5665505160800974
0.9767652237952065   0.4557857901872123   0.7132985675069183   0.2970965932340256   0.6513689084612534   0.8918371870452112   0.49642420383997116   0.8757087070058475   0.3088456066207246   0.8294815523824876   0.9741102119486428   0.43692176757783996   0.14125437653545692   0.8808624177309897   0.915096795260071   0.473053747461687   0.4475033193136792   0.13879435315495706   0.642980558203757   0.7526656828801397   0.568081614696683   0.7690570122313467   0.8891827272104864   0.18611516680004225   0.5913163909014764   0.3132712220441344   0.17588415970356805   0.8890185735660167   0.9399474824402231   0.42143403499892323   0.6794599558635969   0.013309866560169211   0.6311018758194985   0.5919524826164357   0.7053497439149541   0.5763880989823292   0.48984749928404153   0.711090064885446   0.790252948654883   0.10333435152064224   0.04234417997036235   0.5722957117304889   0.14727239045112608   0.3506686686405025   0.47426256527367944   0.8032386994991422   0.25808966324063964   0.16455350184046025   0.8829461743722031   0.4899674774550078   0.08220550353707162   0.2755349282744436   0.94299869193198   0.06853344245608453   0.4027455476734747   0.2622250617142744   0.31189681611248155   0.4765809598396488   0.6973958037585206   0.6858369627319452   0.82204931682844   0.7654908949542029   0.9071428551036375   0.5825026112113029
0.7797051368580776   0.19319518322371396   0.7598704646525114   0.2318339425708004   0.3054425715843982   0.38995648372457176   0.5017808014118718   0.06728044073034015   0.4224963972121951   0.899989006269564   0.41957529787480013   0.7917455124558965   0.47949770528021507   0.8314555638134794   0.016829750201325436   0.5295204507416221   0.16760088916773352   0.35487460397383064   0.3194339464428048   0.843683488009677   0.3455515723392935   0.5893837090196278   0.4122910913391673   0.2611808767983741   0.5658464354812159   0.3961885257959138   0.6524206266866559   0.02934693422757372   0.2604038638968177   0.006232042071342044   0.15063982527478414   0.9620664934972336   0.8379074666846226   0.10624303580177805   0.731064527399984   0.17032098104133703   0.3584097614044075   0.2747874719882986   0.7142347771986586   0.6408005302997148   0.190808872236674   0.9199128680144679   0.3948008307558537   0.7971170422900379   0.8452572998973804   0.3305291589948402   0.9825097394166864   0.5359361654916638   0.2794108644161646   0.9343406331989264   0.3300891127300305   0.5065892312640901   0.019007000519346867   0.9281085911275844   0.17944928745524635   0.5445227377668564   0.18109953383472427   0.8218655553258063   0.44838476005526234   0.3742017567255194   0.8226897724303167   0.5470780833375077   0.7341499828566038   0.7334012264258045
0.6318809001936427   0.6271652153230397   0.3393491521007501   0.9362841841357666   0.7866236002962623   0.2966360563281995   0.3568394126840637   0.40034801864410297   0.5072127358800977   0.36229542312927315   0.02675029995403323   0.8937587873800129   0.48820573536075085   0.4341868320016888   0.8473010124987869   0.34923604961315646   0.3071062015260266   0.6123212766758825   0.3989162524435245   0.9750342928876371   0.4844164290957098   0.06524319333837479   0.6647662695869208   0.24163306646183252   0.8525355289020671   0.43807797801533505   0.32541711748617064   0.30534888232606583   0.06591192860580478   0.1414419216871355   0.9685777048021069   0.9050008636819629   0.558699192725707   0.7791464985578624   0.9418274048480737   0.011242076301949951   0.07049345736495619   0.3449596665561736   0.0945263923492868   0.6620060266887935   0.7633872558389296   0.7326383898802912   0.6956101399057623   0.6869717338011564   0.27897082674321977   0.6673951965419164   0.030843870318841567   0.44533866733932387   0.4264352978411527   0.2293172185265813   0.705426752832671   0.13998978501325804   0.3605233692353479   0.08787529683944575   0.7368490480305641   0.23498892133129515   0.8018241765096409   0.30872879828158334   0.7950216431824904   0.22374684502934522   0.7313307191446846   0.9637691317254098   0.7004952508332036   0.5617408183405518
0.9679434633057551   0.23113074184511864   0.00488511092744132   0.8747690845393954   0.6889726365625354   0.5637355453032022   0.9740412406085998   0.42943041720007147   0.26253733872138263   0.33441832677662103   0.2686144877759288   0.28944063218681343   0.9020139694860347   0.24654302993717525   0.5317654397453647   0.05445171085551828   0.10018979297639391   0.9378142316555919   0.7367437965628744   0.8307048658261731   0.36885907383170924   0.9740450999301822   0.03624854572967077   0.2689640474856213   0.40091561052595415   0.7429143580850635   0.03136343480222945   0.39419496294622597   0.7119429739634189   0.1791788127818612   0.057322194193629696   0.9647645457461546   0.4494056352420362   0.8447604860052402   0.7887077064177009   0.6753239135593411   0.5473916657560014   0.598217456068065   0.25694226667233616   0.6208722027038228   0.44720187277960755   0.660403224412473   0.5201984701094617   0.7901673368776497   0.07834279894789828   0.6863581244822909   0.483949924379791   0.5212032893920284   0.6774271884219442   0.9434437663972274   0.4525864895775616   0.1270083264458024   0.9654842144585253   0.7642649536153662   0.3952642953839319   0.1622437806996479   0.516078579216489   0.9195044676101259   0.606556588966231   0.48691986714030683   0.9686869134604876   0.3212870115420611   0.34961432229389483   0.8660476644364841
0.5214850406808801   0.6608837871295881   0.829415852184433   0.07588032755883432   0.44314224173298183   0.9745256626472971   0.345465927804642   0.5546770381668059   0.7657150533110377   0.031081896250069737   0.8928794382270805   0.42766871172100357   0.8002308388525124   0.26681694263470357   0.49761514284314856   0.26542493102135567   0.28415225963602336   0.34731247502457757   0.8910585538769176   0.7785050638810488   0.31546534617553573   0.026025463482516494   0.5414442315830228   0.9124573994445648   0.7939803054946556   0.3651416763529285   0.7120283793985898   0.8365770718857305   0.35083806376167376   0.3906160137056313   0.36656245159394774   0.2819000337189245   0.585123010450636   0.3595341174555616   0.4736830133668673   0.854231321997921   0.7848921715981235   0.09271717482085805   0.9760678705237187   0.5888063909765653   0.5007399119621002   0.7454046997962804   0.08500931664680111   0.8103013270955165   0.18527456578656443   0.719379236313764   0.5435650850637783   0.8978439276509517   0.39129426029190884   0.3542375599608355   0.8315367056651886   0.06126685576522122   0.0404561965302351   0.9636215462552041   0.4649742540712408   0.7793668220462967   0.4553331860795991   0.6040874287996426   0.9912912407043736   0.9251355000483757   0.6704410144814755   0.5113702539787846   0.015223370180654828   0.3363291090718104
0.1697011025193754   0.765965554182504   0.9302140535338537   0.526027781976294   0.984426536732811   0.046586317868740054   0.3866489684700754   0.6281838543253423   0.5931322764409022   0.6923487579079045   0.5551122628048868   0.566916998560121   0.552676079910667   0.7287272116527004   0.09013800873364596   0.7875501765138243   0.09734289383106792   0.12463978285305775   0.09884676802927242   0.8624146764654486   0.4269018793495924   0.6132695288742732   0.08362339784861758   0.5260855673936382   0.25720077683021697   0.8473039746917692   0.15340934431476388   0.00005778541734421938   0.27277424009740603   0.8007176568230291   0.7667603758446885   0.37187393109200195   0.679641963656504   0.10836889891512459   0.2116481130398017   0.8049569325318809   0.12696588374583692   0.37964168726242425   0.12151010430615573   0.01740675601805654   0.029622989914768992   0.2550019044093665   0.022663336276883314   0.15499207955260794   0.6027211105651766   0.6417323755350932   0.9390399384282657   0.6289065121589698   0.3455203337349596   0.7944284008433241   0.7856305941135019   0.6288487267416255   0.07274609363755358   0.993710744020295   0.018870218268813365   0.2569747956496236   0.39310412998104965   0.8853418451051703   0.8072221052290117   0.4520178631177427   0.2661382462352127   0.5057001578427461   0.6857120009228559   0.43461110709968614
0.23651525632044373   0.25069825343337965   0.6630486646459727   0.27961902754707824   0.6337941457552672   0.6089658778982864   0.7240087262177068   0.6507125153881085   0.2882738120203075   0.8145374770549623   0.9383781321042051   0.021863788646482932   0.21552771838275392   0.8208267330346674   0.9195079138353917   0.7648889929968593   0.8224235884017043   0.9354848879294969   0.11228580860638   0.31287112987911664   0.5562853421664915   0.42978473008675083   0.42657380768352404   0.8782600227794305   0.3197700858460478   0.17908647665337116   0.7635251430375515   0.5986409952323523   0.6859759400907807   0.5701205987550848   0.03951641681984454   0.9479284798442438   0.39770212807047317   0.7555831217001224   0.10113828471563949   0.9260646911977608   0.18217440968771925   0.9347563886654551   0.1816303708802478   0.16117569820090152   0.359750821286015   0.9992715007359582   0.0693445622738678   0.8483045683217849   0.8034654791195234   0.5694867706492074   0.6427707545903437   0.9700445455423544   0.4836953932734756   0.3904002939958362   0.8792456115527923   0.3714035503100021   0.7977194531826949   0.8202796952407514   0.8397291947329478   0.42347507046575833   0.40001732511222177   0.06469657354062898   0.7385909100173083   0.49741037926799747   0.2178429154245025   0.12994018487517386   0.5569605391370605   0.336234681067096
0.8580920941384875   0.1306686841392157   0.48761597686319264   0.4879301127453111   0.054626615018964084   0.5611819134900083   0.8448452222728489   0.5178855672029568   0.5709312217454885   0.17078161949417217   0.9655996107200566   0.1464820168929546   0.7732117685627935   0.35050192425342075   0.12587041598710882   0.7230069464271962   0.3731944434505718   0.2858053507127918   0.38727950596980054   0.22559656715919876   0.1553515280260693   0.15586516583761792   0.8303189668327401   0.8893618860921028   0.2972594338875818   0.02519648169840221   0.34270298996954746   0.4014317733467917   0.2426328188686177   0.4640145682083938   0.49785776769669854   0.883546206143835   0.6717015971231293   0.2932329487142217   0.5322581569766419   0.7370641892508804   0.8984898285603357   0.9427310244608009   0.40638774098953306   0.01405724282368416   0.5252953851097639   0.6569256737480091   0.01910823501973252   0.7884606756644854   0.3699438570836946   0.5010605079103913   0.18878926818699243   0.8990987895723827   0.0726844231961128   0.475864026211989   0.846086278217445   0.49766701622559095   0.8300516043274951   0.01184945800359514   0.3482285105207465   0.614120810081756   0.15835000720436587   0.7186165092893735   0.8159703535441045   0.8770566208308755   0.25986017864403016   0.7758854848285726   0.40958261255457146   0.8629993780071914
0.7345647935342663   0.11895981108056346   0.39047437753483893   0.074538702342706   0.3646209364505717   0.6178993031701723   0.20168510934784653   0.17543991277032336   0.29193651325445885   0.14203527695818327   0.3555988311304015   0.6777728965447324   0.46188490892696377   0.13018581895458814   0.007370320609655073   0.06365208646297646   0.3035349017225979   0.41156930966521466   0.1913999670655505   0.1865954656321009   0.04367472307856771   0.6356838248366421   0.781817354510979   0.3235960876249095   0.30910992954430144   0.5167240137560786   0.39134297697614007   0.2490573852822035   0.9444889930937298   0.8988247105859064   0.18965786762829356   0.07361747251188012   0.6525524798392709   0.7567894336277231   0.834059036497892   0.39584457596714767   0.19066757091230713   0.626603614673135   0.8266887158882369   0.33219248950417124   0.8871326691897092   0.21503430500792028   0.6352887488226864   0.14559702387207032   0.8434579461111416   0.5793504801712782   0.8534713943117074   0.8220009362471609   0.5343480165668401   0.0626264664151996   0.4621284173355673   0.5729435509649573   0.5898590234731104   0.16380175582929324   0.27247054970727375   0.49932607845307725   0.9373065436338395   0.40701232220157013   0.4384115132093817   0.10348150248592954   0.7466389727215322   0.7804087075284352   0.6117227973211448   0.7712890129817583
0.859506303531823   0.565374402520515   0.9764340484984584   0.6256919891096879   0.016048357420681503   0.9860239223492366   0.12296265418675098   0.8036910528625272   0.4817003408538414   0.9233974559340371   0.6608342368511837   0.2307475018975698   0.8918413173807311   0.7595957001047439   0.38836368714390995   0.7314214234444926   0.9545347737468917   0.3525833779031737   0.9499521739345282   0.627939920958563   0.2078958010253594   0.5721746703747385   0.3382293766133834   0.8566509079768048   0.34838949749353637   0.006800267854223593   0.36179532811492504   0.23095891886711675   0.33234114007285487   0.0207763455049869   0.2388326739281741   0.4272678660045896   0.8506407992190135   0.09737888957094981   0.5779984370769904   0.19652036410701978   0.9587994818382823   0.33778318946620595   0.18963474993308044   0.4650989406625272   0.004264708091390672   0.9851998115630323   0.23968257599855222   0.8371590197039642   0.7963689070660313   0.41302514118829375   0.9014531993851688   0.9805081117271595   0.44797940957249494   0.40622487333407015   0.5396578712702438   0.7495491928600427   0.11563826949964007   0.38544852782908323   0.30082519734206964   0.32228132685545313   0.26499747028062665   0.2880696382581334   0.7228267602650793   0.12576096274843332   0.30619798844234425   0.9502864487919275   0.5331920103319988   0.6606620220859061
0.3019332803509536   0.9650866372288952   0.29350943433344656   0.823503002381942   0.5055643732849223   0.5520614960406015   0.3920562349482778   0.8429948906547825   0.057584963712427405   0.14583662270653133   0.852398363678034   0.09344569779473973   0.9419466942127873   0.7603880948774481   0.5515731663359644   0.7711643709392866   0.6769492239321607   0.47231845661931465   0.8287464060708851   0.6454034081908533   0.3707512354898165   0.5220320078273871   0.2955543957388863   0.9847413861049472   0.06881795513886285   0.5569453705984919   0.0020449614054397335   0.16123838372300525   0.5632535818539405   0.00488387455789042   0.609988726457162   0.3182434930682228   0.5056686181415131   0.8590472518513591   0.757590362779128   0.22479779527348306   0.5637219239287258   0.09865915697391099   0.20601719644316352   0.45363342433419646   0.886772699996565   0.6263407003545963   0.3772707903722784   0.8082300161433432   0.5160214645067486   0.10430869252720917   0.08171639463339207   0.823488630038396   0.4472035093678858   0.5473633219287173   0.07967143322795234   0.6622502463153908   0.8839499275139452   0.5424794473708269   0.4696827067707904   0.344006753247168   0.3782813093724321   0.6834321955194678   0.7120923439916624   0.11920895797368494   0.8145593854437063   0.5847730385455567   0.5060751475484989   0.6655755336394885
0.9277866854471413   0.9584323381909604   0.12880435717622057   0.8573455174961453   0.4117652209403927   0.8541236456637513   0.0470879625428285   0.03385688745774923   0.9645617115725069   0.30676032373503404   0.9674165293148762   0.3716066411423584   0.08061178405856169   0.7642808763642072   0.49773382254408577   0.027599887895190422   0.7023304746861296   0.08084868084473941   0.7856414785524233   0.9083909299215055   0.8877710892424232   0.49607564229918266   0.2795663310039243   0.242815396282017   0.9599844037952819   0.5376433041082221   0.15076197382770376   0.38546987878587174   0.5482191828548894   0.6835196584444709   0.10367401128487526   0.3516129913281225   0.5836574712823824   0.3767593347094369   0.1362574819699991   0.9800063501857641   0.5030456872238207   0.6124784583452297   0.6385236594259133   0.9524064622905737   0.8007152125376911   0.5316297775004903   0.85288218087349   0.04401553236906818   0.9129441232952679   0.0355541352013077   0.5733158498695657   0.8012001360870512   0.9529597194999858   0.49791083109308554   0.42255387604186195   0.4157302573011794   0.40474053664509657   0.8143911726486146   0.3188798647569867   0.0641172659730569   0.8210830653627141   0.43763183793917765   0.18262238278698759   0.08411091578729282   0.3180373781388935   0.825153379593948   0.5440987233610742   0.13170445349671916
0.5173221656012024   0.29352360209345757   0.6912165424875842   0.08768892112765098   0.6043780423059345   0.2579694668921499   0.11790069261801853   0.2864887850405998   0.6514183228059487   0.7600586357990644   0.6953468165761566   0.8707585277394204   0.24667778616085215   0.9456674631504498   0.3764669518191699   0.8066412617663634   0.425594720798138   0.5080356252112721   0.1938445690321823   0.7225303459790706   0.10755734265924448   0.6828822456173242   0.649745845671108   0.5908258924823515   0.5902351770580421   0.3893586435238666   0.9585293031835238   0.5031369713547005   0.9858571347521076   0.13138917663171676   0.8406286105655053   0.2166481863141007   0.3344388119461588   0.3713305408326524   0.14528179398934868   0.34588965857468035   0.0877610257853067   0.42566307768220263   0.7688148421701788   0.5392483968083169   0.6621663049871688   0.9176274524709305   0.5749702731379965   0.8167180508292462   0.5546089623279242   0.2347452068536063   0.9252244274668885   0.22589215834689477   0.9643737852698822   0.8453865633297397   0.9666951242833647   0.7227551869921942   0.9785166505177746   0.7139973866980229   0.12606651371785935   0.5061070006780936   0.6440778385716158   0.3426668458653705   0.9807847197285107   0.1602173421034132   0.5563168127863091   0.9170037681831679   0.21196987755833188   0.6209689452950963
0.8941505077991404   0.9993763157122374   0.6369996044203354   0.8042508944658501   0.3395415454712161   0.7646311088586311   0.7117751769534469   0.5783587361189553   0.3751677602013339   0.9192445455288915   0.7450800526700824   0.8556035491267611   0.39665110968355927   0.20524715883086853   0.619013538952223   0.3494965484486675   0.7525732711119435   0.862580312965498   0.6382288192237123   0.1892792063452543   0.1962564583256344   0.9455765447823301   0.4262589416653804   0.5683102610501579   0.302105950526494   0.9462002290700927   0.789259337245045   0.7640593665843078   0.962564405055278   0.1815691202114616   0.0774841602915981   0.1857006304653526   0.587396644853944   0.26232457468257014   0.3324041076215158   0.33009708133859156   0.19074553517038473   0.05707741585170162   0.7133905686692928   0.980600532889924   0.43817226405844123   0.19449710288620362   0.0751617494455805   0.7913213265446698   0.24191580573280683   0.2489205581038735   0.6489028077802   0.22301106549451177   0.9398098552063128   0.3027203290337808   0.859643470535155   0.4589516989102039   0.9772454501510348   0.1211512088223192   0.7821593102435569   0.2732510684448513   0.3898488052970908   0.858826634139749   0.4497552026220411   0.9431539871062598   0.19910327012670612   0.8017492182880475   0.7363646339527483   0.9625534542163358
0.7609310060682649   0.6072521154018439   0.6612028845071678   0.17123212767166596   0.519015200335458   0.35833155729797034   0.012300076726967736   0.9482210621771542   0.5792053451291452   0.05561122826418952   0.15265660619181273   0.4892693632669503   0.6019598949781104   0.9344600194418703   0.3704972959482558   0.21601829482209903   0.21211108968101955   0.07563338530212127   0.9207420933262147   0.27286430771583925   0.013007819554313427   0.27388416701407386   0.1843774593734664   0.31031085349950355   0.25207681348604855   0.66663205161223   0.5231745748662986   0.1390787258278376   0.7330616131505905   0.3083004943142597   0.5108744981393308   0.1908576636506834   0.1538562680214453   0.2526892660500702   0.35821789194751813   0.7015883003837331   0.5518963730433349   0.31822924660819984   0.9877205959992623   0.4855700055616341   0.3397852833623154   0.24259586130607858   0.06697850267304761   0.21270569784579482   0.32677746380800193   0.9687116942920048   0.8826010432995812   0.9023948443462912   0.0747006503219534   0.3020796426797747   0.35942646843328263   0.7633161185184536   0.34163903717136285   0.9937791483655151   0.8485519702939518   0.5724584548677703   0.18778276914991757   0.7410898823154448   0.49033407834643367   0.8708701544840372   0.6358863961065826   0.42286063570724497   0.5026134823471714   0.38530014892240305
0.29610111274426726   0.1802647744011664   0.43563497967412373   0.1725944510766082   0.9693236489362653   0.21155308010916166   0.5530339363745426   0.27019960673031695   0.8946229986143119   0.9094734374293869   0.19360746794125988   0.5068834882118634   0.552983961442949   0.9156942890638718   0.3450554976473081   0.9344250333440931   0.36520119229303144   0.17460440674842706   0.8547214193008744   0.06355487886005594   0.7293147961864488   0.7517437710411821   0.352107936953703   0.6782547299376529   0.43321368344218153   0.5714789966400157   0.9164729572795792   0.5056602788610447   0.4638900345059162   0.35992591653085404   0.36343902090503677   0.23546067213072772   0.5692670358916043   0.45045247910146713   0.16983155296377686   0.7285771839188644   0.016283074448655302   0.5347581900375952   0.8247760553164688   0.7941521505747714   0.6510818821556239   0.36015378328916814   0.9700546360155944   0.7305972717147154   0.921767085969175   0.6084100122479861   0.6179466990618914   0.05234254177706253   0.48855340252699353   0.0369310156079704   0.7014737417823121   0.5466822629160178   0.024663368021077284   0.6770050990771164   0.33803472087727543   0.3112215907852901   0.45539633212947295   0.22655261997564927   0.16820316791349854   0.5826444068664257   0.43911325768081766   0.6917944299380541   0.34342711259702974   0.7884922562916543
0.7880313755251938   0.33164064664888593   0.3733724765814353   0.05789498457693891   0.8662642895560188   0.7232306344008999   0.7554257775195439   0.005552442799876376   0.3777108870290252   0.6862996187929294   0.053952035737231736   0.45887017988385853   0.35304751900794795   0.009294519715813075   0.7159173148599564   0.1476485890985684   0.897651186878475   0.7827418997401638   0.5477141469464578   0.5650041822321427   0.45853792919765735   0.09094746980210973   0.20428703434942808   0.7765119259404883   0.6705065536724636   0.7593068231532238   0.8309145577679927   0.7186169413635495   0.8042422641164448   0.03607618875232396   0.07548878024844889   0.713064498563673   0.42653137708741956   0.3497765699593945   0.021536744511217152   0.25419431867981457   0.07348385807947161   0.3404820502435814   0.3056194296512608   0.10654572958124615   0.1758326712009966   0.5577401505034176   0.7579052827048031   0.5415415473491034   0.7172947420033393   0.4667926807013079   0.553618248355375   0.7650296214086151   0.04678818833087572   0.7074858575480841   0.7227036905873822   0.0464126800450656   0.2425459242144309   0.6714096687957601   0.6472149103389333   0.3333481814813925   0.8160145471270114   0.3216330988363656   0.6256781658277161   0.07915386280157795   0.7425306890475397   0.9811510485927841   0.3200587361764553   0.9726081332203318
0.5666980178465432   0.42341089808936655   0.5621534534716522   0.4310665858712283   0.8494032758432039   0.9566182173880586   0.008535205116277342   0.6660369644626133   0.8026150875123281   0.24913235983997456   0.28583151452889516   0.6196242844175477   0.5600691632978972   0.5777226910442144   0.6386166041899619   0.28627610293615513   0.7440546161708859   0.25608959220784877   0.012938438362245782   0.20712224013457722   0.0015239271233461473   0.2749385436150646   0.6928797021857904   0.23451410691424543   0.43482590927680304   0.851527645525698   0.13072624871413818   0.8034475210430171   0.5854226334335991   0.8949094281376394   0.12219104359786084   0.13741055658040383   0.782807545921271   0.6457770682976649   0.8363595290689657   0.5177862721628561   0.2227383826233738   0.06805437725345047   0.19774292487900377   0.23151016922670098   0.4786837664524879   0.8119647850456017   0.184804486516758   0.024387929092123783   0.47715983932914174   0.537026241430537   0.4919247843309675   0.7898738221778784   0.04233393005233874   0.685498595904839   0.3611985356168293   0.9864263011348613   0.4569112966187396   0.7905891677671996   0.23900749201896845   0.8490157445544575   0.6741037506974685   0.14481209946953466   0.4026479629500028   0.33122947239160133   0.4513653680740947   0.0767577222160842   0.20490503807099902   0.09971930316490032
0.9726816016216068   0.2647929371704825   0.020100551554241054   0.07533137407277654   0.49552176229246503   0.7277666957399455   0.5281757672232735   0.2854575518948982   0.4531878322401263   0.0422680998351065   0.16697723160644423   0.2990312507600369   0.9962765356213867   0.251678932067907   0.9279697395874758   0.45001550620557945   0.3221727849239182   0.10686683259837229   0.5253217766374729   0.11878603381397812   0.8708074168498234   0.030109110382288085   0.32041673856647396   0.019066730649077795   0.8981258152282167   0.7653161732118056   0.3003161870122329   0.9437353565763013   0.4026040529357516   0.03754947747186007   0.7721404197889593   0.6582778046814031   0.9494162206956253   0.9952813776367536   0.6051631881825151   0.3592465539213662   0.9531396850742385   0.7436024455688466   0.6771934485950394   0.9092310477157868   0.6309669001503203   0.6367356129704743   0.15187167195756637   0.7904450139018087   0.7601594833004969   0.6066265025881863   0.8314549333910924   0.7713782832527308   0.8620336680722802   0.8413103293763807   0.5311387463788595   0.8276429266764296   0.4594296151365287   0.8037608519045206   0.7589983265899002   0.16936512199502649   0.5100133944409034   0.808479474267767   0.1538351384073851   0.8101185680736603   0.5568737093666649   0.06487702869892044   0.4766416898123458   0.9008875203578736
0.9259068092163446   0.4281414157284461   0.3247700178547794   0.11044250645606495   0.1657473259158477   0.8215149131402598   0.493315084463687   0.3390642232033341   0.3037136578435674   0.9802045837638792   0.9621763380848274   0.5114212965269046   0.8442840427070387   0.17644373185935858   0.20317801149492723   0.3420561745318781   0.33427064826613534   0.3679642575915915   0.04934287308754215   0.5319376064582177   0.7773969388994704   0.3030872288926711   0.5727011832751964   0.6310500861003442   0.8514901296831259   0.8749458131642249   0.247931165420417   0.5206075796442793   0.6857428037672781   0.0534309000239651   0.75461608095673   0.1815433564409451   0.3820291459237107   0.07322631626008591   0.7924397428719026   0.6701220599140405   0.5377451032166719   0.8967825844007273   0.5892617313769754   0.32806588538216247   0.20347445495053662   0.5288183268091359   0.5399188582894332   0.7961282789239447   0.42607751605106625   0.22573109791646476   0.9672176750142368   0.16507819282360053   0.5745873863679404   0.3507852847522398   0.7192865095938198   0.6444706131793213   0.8888445826006622   0.2973543847282747   0.9646704286370898   0.4629272567383762   0.5068154366769516   0.22412806846818878   0.1722306857651872   0.7928051968243357   0.9690703334602796   0.32734548406746145   0.582968954388212   0.4647393114421732
0.765595878509743   0.7985271572583256   0.04305009609877872   0.6686110325182285   0.3395183624586768   0.5727960593418608   0.07583242108454193   0.5035328396946279   0.7649309760907363   0.22201077458962104   0.3565459114907221   0.8590622265153066   0.8760863934900741   0.9246563898613464   0.39187548285363233   0.3961349697769304   0.3692709568131225   0.7005283213931576   0.2196447970884451   0.6033297729525947   0.40020062335284284   0.3731828373256961   0.6366758427002333   0.13859046151042156   0.6346047448430998   0.5746556800673706   0.5936257466014545   0.4699794289921931   0.2950863823844231   0.0018596207255097248   0.5177933255169126   0.9664465892975652   0.5301554062936867   0.7798488461358887   0.16124741402619044   0.10738436278225855   0.6540690128036126   0.8551924562745423   0.7693719311725581   0.7112493930053282   0.28479805599049013   0.15466413488138475   0.549727134084113   0.1079196200527334   0.8845974326376472   0.7814812975556886   0.9130512913838799   0.9693291585423118   0.24999268779454742   0.20682561748831804   0.31942554478242535   0.49934972955011875   0.9549063054101243   0.20496599676280833   0.8016322192655128   0.5329031402525536   0.42475089911643765   0.4251171506269196   0.6403848052393223   0.425518777470295   0.7706818863128251   0.5699246943523774   0.8710128740667642   0.7142693844649669
0.4858838303223349   0.41526055947099255   0.32128573998265114   0.6063497644122334   0.6012863976846876   0.633779261915304   0.40823444859877134   0.6370206058699216   0.35129370989014025   0.4269536444269859   0.08880890381634599   0.13767087631980293   0.3963874044800159   0.22198764766417758   0.28717668455083323   0.6047677360672493   0.9716365053635783   0.796870497037258   0.6467918793115108   0.17924895859695436   0.20095461905075326   0.22694580268488065   0.7757790052447467   0.4649795741319875   0.7150707887284183   0.8116852432138881   0.45449326526209555   0.858629809719754   0.11378439104373067   0.17790598129858412   0.04625881666332421   0.22160920384983238   0.7624906811535904   0.7509523368715982   0.9574499128469782   0.08393832753002944   0.3661032766735745   0.5289646892074206   0.670273228296145   0.47917059146278007   0.3944667713099962   0.7320941921701627   0.02348134898463413   0.29992163286582574   0.19351215225924295   0.5051483894852821   0.24770234373988745   0.8349420587338382   0.4784413635308246   0.6934631462713939   0.7932090784777919   0.9763122490140842   0.36465697248709394   0.5155571649728098   0.7469502618144677   0.7547030451642519   0.6021662913335035   0.7646048281012116   0.7895003489674894   0.6707647176342224   0.23606301465992904   0.23564013889379098   0.11922712067134446   0.19159412617144234
0.8415962433499329   0.5035459467236283   0.09574577168671032   0.8916724933056166   0.6480840910906899   0.9983975572383462   0.8480434279468229   0.056730434571778364   0.16964272755986531   0.30493441096695234   0.05483434946903098   0.08041818555769413   0.8049857550727714   0.7893772459941425   0.30788408765456327   0.32571514039344224   0.20281946373926785   0.024772417892930925   0.5183837386870738   0.6549504227592198   0.9667564490793388   0.78913227899914   0.3991566180157293   0.4633562965877775   0.12516020572940595   0.28558633227551167   0.30341084632901905   0.5716838032821608   0.477076114638716   0.2871887750371654   0.45536741838219613   0.5149533687103826   0.3074333870788507   0.982254364070213   0.40053306891316515   0.43453518315268835   0.5024476320060793   0.19287711807607053   0.09264898125860188   0.10882004275924612   0.2996281682668115   0.16810470018313958   0.5742652425715281   0.4538696200000263   0.3328717191874727   0.37897242118399965   0.1751086245557987   0.9905133234122488   0.20771151345806677   0.09338608890848799   0.8716977782267797   0.41882952013008795   0.7306353988193508   0.8061973138713227   0.41633035984458355   0.9038761514197055   0.42320201174050004   0.8239429498011096   0.015797290931418385   0.4693409682670171   0.9207543797344208   0.631065831725039   0.9231483096728165   0.360520925507771
0.6211262114676093   0.4629611315418995   0.34888306710128847   0.9066513055077446   0.2882544922801365   0.08398871035789984   0.17377444254548974   0.9161379820954959   0.08054297882206975   0.9906026214494118   0.30207666431871005   0.4973084619654079   0.349907580002719   0.18440530757808923   0.8857463044741265   0.5934323105457024   0.926705568262219   0.36046235777697966   0.8699490135427081   0.12409134227868539   0.005951188527798254   0.7293965260519406   0.9468007038698916   0.7635704167709144   0.38482497706018903   0.2664353945100411   0.5979176367686032   0.8569191112631698   0.09657048478005253   0.18244668415214124   0.4241431942231134   0.9407811291676739   0.016027505957982784   0.1918440627027294   0.12206652990440339   0.44347266720226597   0.6661199259552638   0.007438755124640176   0.2363202254302769   0.8500403566565635   0.7394143576930449   0.6469763973476605   0.36637121188756877   0.7259490143778782   0.7334631691652466   0.9175798712957199   0.41957050801767715   0.9623785976069636   0.34863819210505753   0.6511444767856789   0.821652871249074   0.10545948634379394   0.252067707325005   0.4686977926335376   0.3975096770259606   0.16467835717612006   0.23604020136702222   0.2768537299308082   0.2754431471215572   0.721205689973854   0.5699202754117584   0.26941497480616805   0.0391229216912803   0.8711653333172905
0.8305059177187136   0.6224385774585075   0.6727517098037116   0.14521631893941242   0.09704274855346703   0.7048587061627876   0.25318120178603437   0.18283772133244874   0.7484045564484095   0.05371422937710867   0.4315283305369603   0.07737823498865479   0.49633684912340453   0.5850164367435711   0.03401865351099975   0.9126998778125347   0.2602966477563823   0.30816270681276287   0.7585755063894426   0.19149418783868066   0.6903763723446239   0.03874773200659481   0.7194525846981623   0.3203288545213901   0.8598704546259103   0.4163091545480873   0.04670087489445074   0.17511253558197767   0.7628277060724432   0.7114504483852998   0.7935196731084164   0.9922748142495289   0.014423149624033705   0.6577362190081911   0.36199134257145604   0.9148965792608742   0.5180863005006292   0.07271978226462003   0.3279726890604563   0.0021967014483394148   0.2577896527442469   0.7645570754518571   0.5693971826710137   0.8107025136096587   0.567413280399623   0.7258093434452624   0.8499445979728515   0.49037365908826863   0.7075428257737127   0.30950018889717507   0.8032437230784008   0.315261123506291   0.9447151197012695   0.5980497405118753   0.009724049969984343   0.3229863092567621   0.9302919700772359   0.9403135215036842   0.6477327073985283   0.40808972999588794   0.4122056695766067   0.8675937392390642   0.319760018338072   0.4058930285475485
0.15441601683235978   0.10303666378720701   0.7503628356670582   0.5951905149378898   0.5870027364327367   0.3772273203419446   0.9004182376942068   0.10481685584962108   0.879459910659024   0.06772713144476955   0.09717451461580603   0.7895557323433301   0.9347447909577543   0.46967739093289423   0.0874504646458217   0.466569423086568   0.004452820880518481   0.52936386942921   0.4397177572472934   0.05847969309068011   0.5922471513039118   0.6617701301901457   0.11995773890922141   0.6525866645431316   0.43783113447155203   0.5587334664029387   0.36959490324216315   0.057396149605241864   0.8508283980388153   0.18150614606099413   0.4691766655479564   0.9525792937556208   0.9713684873797913   0.1137790146162246   0.3720021509321504   0.16302356141229069   0.036623696422037014   0.6441016236833303   0.28455168628632865   0.6964541383257227   0.03217087554151853   0.11473775425412037   0.8448339290390353   0.6379744452350425   0.43992372423760673   0.45296762406397456   0.7248761901298139   0.9853877806919109   0.0020925897660546973   0.8942341576610358   0.35528128688765065   0.927991631086669   0.1512641917272394   0.7127280116000416   0.8861046213396943   0.9754123373310483   0.17989570434744803   0.5989489969838171   0.5141024704075439   0.8123887759187576   0.143272007925411   0.9548473733004867   0.22955078412121524   0.11593463759303495
0.11110113238389248   0.8401096190463663   0.38471685508217995   0.4779601923579924   0.6711774081462858   0.38714199498239177   0.6598406649523662   0.49257241166608146   0.669084818380231   0.49290783732135596   0.30455937806471545   0.5645807805794124   0.5178206266529917   0.7801798257213143   0.4184547567250212   0.589168443248364   0.33792492230554366   0.1812308287374972   0.9043522863174772   0.7767796673296065   0.19465291438013263   0.22638345543701052   0.674801502196262   0.6608450297365716   0.08355178199624014   0.38627383639064417   0.29008464711408205   0.18288483737857913   0.4123743738499544   0.9991318414082524   0.630243982161716   0.6903124257124977   0.7432895554697233   0.5062240040868965   0.3256846040970005   0.1257316451330853   0.22546892881673167   0.7260441783655822   0.9072298473719793   0.5365632018847212   0.887544006511188   0.544813349628085   0.00287756105450206   0.7597835345551147   0.6928910921310554   0.31842989419107454   0.32807605885824004   0.09893850481854322   0.6093393101348152   0.9321560578004303   0.03799141174415799   0.9160536674399641   0.1969649362848609   0.9330242163921779   0.40774742958244203   0.2257412417274664   0.4536753808151376   0.42680021230528137   0.08206282548544157   0.10000959659438109   0.22820645199840592   0.7007560339396991   0.17483297811346224   0.5634463947096598
0.3406624454872179   0.15594268431161412   0.1719554170589602   0.8036628601545451   0.6477713533561625   0.8375127901205396   0.8438793582007201   0.704724355336002   0.038432043221347224   0.9053567323201093   0.8058879464565621   0.7886706878960379   0.8414671069364863   0.9723325159279314   0.3981405168741201   0.5629294461685714   0.38779172612134877   0.54553230362265   0.31607769138867853   0.46291984957419036   0.15958527412294288   0.8447762696829508   0.1412447132752163   0.8994734548645305   0.818922828635725   0.6888335853713368   0.9692892962162561   0.09581059470998535   0.17115147527956248   0.8513207952507972   0.12540993801553593   0.3910862393739834   0.13271943205821526   0.9459640629306879   0.31952199155897376   0.6024155514779456   0.29125232512172894   0.9736315470027566   0.9213814746848537   0.03948610530937413   0.9034605990003801   0.4280992433801065   0.6053037832961752   0.5765662557351837   0.7438753248774372   0.5833229736971557   0.46405907002095886   0.6770928008706533   0.9249524962417123   0.8944893883258189   0.4947697738047027   0.581282206160668   0.7538010209621498   0.04316859307502179   0.3693598357891668   0.19019596678668452   0.6210815889039345   0.0972045301443339   0.049837844230193024   0.5877804153087389   0.3298292637822056   0.12357298314157739   0.12845636954533934   0.5482943099993648
0.42636866478182545   0.6954737397614709   0.5231525862491643   0.9717280542641811   0.6824933399043882   0.11215076606431516   0.05909351622820539   0.29463525339352775   0.7575408436626759   0.21766137773849623   0.5643237424235027   0.7133530472328599   0.003739822700526071   0.17449278466347443   0.19496390663433585   0.5231570804461753   0.38265823379659153   0.07728825451914052   0.14512606240414283   0.9353766651374363   0.052828970014385905   0.9537152713775632   0.016669692858803466   0.3870823551380716   0.6264603052325605   0.2582415316160923   0.4935171066096392   0.4153543008738906   0.9439669653281723   0.14609076555177714   0.43442359038143386   0.12071904748036283   0.18642612166549638   0.9284293878132809   0.8700998479579312   0.407366000247503   0.1826862989649703   0.7539366031498065   0.6751359413235953   0.8842089198013278   0.8000280651683788   0.6766483486306659   0.5300098789194525   0.9488322546638913   0.7471990951539929   0.7229330772531029   0.5133401860606491   0.5617498995258198   0.12073878992143243   0.46469154563701054   0.019823079451009838   0.1463955986519292   0.17677182459326016   0.3186007800852334   0.585399489069576   0.025676551171566368   0.9903457029277638   0.3901713922719525   0.7152996411116448   0.6183105509240634   0.8076594039627935   0.636234789122146   0.04016369978804942   0.7341016311227356
0.007631338794414722   0.95958644049148   0.5101538208685968   0.7852693764588443   0.26043224364042183   0.2366533632383772   0.9968136348079478   0.22351947693302454   0.13969345371898942   0.7719618176013666   0.976990555356938   0.07712387828109535   0.9629216291257292   0.45336103751613327   0.39159106628736196   0.051447327109528984   0.9725759261979655   0.06318964524418076   0.6762914251757172   0.43313677618546564   0.16491652223517198   0.42695485612203476   0.6361277253876678   0.69903514506273   0.15728518344075723   0.4673684156305547   0.1259739045190709   0.9137657686038857   0.8968529398003354   0.2307150523921775   0.12916026971112307   0.6902462916708612   0.757159486081346   0.4587532347908108   0.1521697143541851   0.6131224133897658   0.7942378569556167   0.005392197274677558   0.7605786480668232   0.5616750862802369   0.8216619307576513   0.9422025520304969   0.08428722289110593   0.1285383100947712   0.6567454085224793   0.5152476959084621   0.44815949750343814   0.4295031650320412   0.49946022508172205   0.04787928027790736   0.3221855929843673   0.5157373964281555   0.6026072852813866   0.8171642278857298   0.1930253232732442   0.8254911047572944   0.8454477992000407   0.35841099309491903   0.04085560891905909   0.2123686913675285   0.051209942244423996   0.3530187958202415   0.28027696085223597   0.6506936050872917
0.22954801148677276   0.4108162437897447   0.19598973796113003   0.5221552949925204   0.5728026029642935   0.8955685478812826   0.7478302404576919   0.09265212996047927   0.07334237788257145   0.8476892676033753   0.4256446474733246   0.5769147335323238   0.4707350926011848   0.03052503971764541   0.23261932420008039   0.7514236287750294   0.6252872934011441   0.6721140466227263   0.1917637152810213   0.5390549374075009   0.5740773511567201   0.31909525080248485   0.9114867544287854   0.8883613323202093   0.34452933966994737   0.9082790070127402   0.7154970164676553   0.3662060373276888   0.7717267367056538   0.01271045913145754   0.9676667760099634   0.2735539073672095   0.6983843588230825   0.16502119152808226   0.5420221285366389   0.6966391738348857   0.22764926622189763   0.13449615181043686   0.3094028043365585   0.9452155450598563   0.6023619728207535   0.4623821051877105   0.11763908905553719   0.4061606076523554   0.028284621664033414   0.14328685438522562   0.20615233462675184   0.5177992753321461   0.6837552819940861   0.23500784737248545   0.4906553181590965   0.15159323800445734   0.9120285452884321   0.2222973882410279   0.522988542149133   0.8780393306372478   0.21364418646534974   0.05727619671294565   0.9809664136124941   0.18140015680236207   0.9859949202434521   0.9227800449025088   0.6715636092759357   0.23618461174250577
0.3836329474226986   0.4603979397147983   0.5539245202203985   0.8300240040901504   0.3553483257586652   0.31711108532957266   0.34777218559364664   0.3122247287580043   0.6715930437645791   0.08210323795708722   0.8571168674345501   0.16063149075354693   0.7595644984761469   0.8598058497160593   0.3341283252854171   0.2825921601162991   0.5459203120107972   0.8025296530031136   0.3531619116729229   0.10119200331393706   0.559925391767345   0.8797496081006049   0.6815983023969873   0.8650073915714313   0.17629244434464647   0.41935166838580656   0.12767378217658873   0.0349833874812809   0.8209441185859813   0.10224058305623389   0.7799015965829421   0.7227586587232766   0.14935107482140217   0.020137345099146654   0.9227847291483919   0.5621271679697297   0.3897865763452552   0.16033149538308733   0.5886564038629749   0.27953500785343055   0.843866264334458   0.3578018423799737   0.235494492190052   0.1783430045394935   0.283940872567113   0.4780522342793688   0.5538961897930648   0.3133356129680622   0.10764842822246651   0.05870056589356224   0.42622240761647606   0.2783522254867813   0.28670430963648524   0.9564599828373284   0.646320811033534   0.5555935667635047   0.13735323481508308   0.9363226377381817   0.723536081885142   0.993466398793775   0.7475666584698278   0.7759911423550944   0.13487967802216705   0.7139313909403444
0.9037003941353698   0.4181892999751207   0.899385185832115   0.5355883864008509   0.6197595215682569   0.9401370656957518   0.34548899603905026   0.2222527734327887   0.5121110933457903   0.8814364998021896   0.9192665884225742   0.9439005479460074   0.2254067837093051   0.9249765169648613   0.27294577738904024   0.38830698118250273   0.08805354889422201   0.9886538792266796   0.5494096955038983   0.3948405823887277   0.3404868904243942   0.2126627368715852   0.41453001748173124   0.6809091914483832   0.4367864962890244   0.7944734368964645   0.5151448316496162   0.1453208050475324   0.8170269747207676   0.8543363712007126   0.16965583561056594   0.9230680316147437   0.3049158813749772   0.972899871398523   0.2503892471879917   0.9791674836687363   0.07950909766567214   0.04792335443366169   0.9774434697989515   0.5908605024862336   0.9914555487714501   0.059269475206982114   0.4280337742950532   0.19601992009750588   0.650968658347056   0.8466067383353969   0.01350375681332198   0.5151107286491226   0.2141821620580316   0.0521333014389324   0.4983589251637058   0.3697899236015902   0.39715518733726407   0.1977969302382198   0.32870308955313987   0.44672189198684653   0.09223930596228681   0.2248970588396968   0.07831384236514816   0.4675544083181102   0.012730208296614668   0.1769737044060351   0.10087037256619667   0.8766939058318766
0.021274659525164538   0.11770422919905299   0.6728365982711435   0.6806739857343708   0.3703060011781086   0.2710974908636561   0.6593328414578215   0.16556325708524813   0.156123839120077   0.21896418942472368   0.1609739162941157   0.795773333483658   0.7589686517828129   0.021167259186503907   0.8322708267409759   0.34905144149681144   0.6667293458205261   0.7962702003468071   0.7539569843758277   0.8814970331787012   0.6539991375239115   0.619296495940772   0.653086611809631   0.004803127346824632   0.632724477998747   0.501592266741719   0.9802500135384875   0.32412914161245393   0.26241847682063835   0.2304947758780629   0.320917172080666   0.15856588452720577   0.10629463770056136   0.01153058645333924   0.1599432557865503   0.36279255104354785   0.3473259859177484   0.9903633272668353   0.3276724290455745   0.013741109546736406   0.6805966400972222   0.19409312692002822   0.5737154446697468   0.13224407636803517   0.026597502573310783   0.5747966309792563   0.9206288328601159   0.12744094902121053   0.39387302457456386   0.07320436423753722   0.9403788193216284   0.8033118074087566   0.1314545477539255   0.8427095883594743   0.6194616472409623   0.6447459228815509   0.02515991005336415   0.831179001906135   0.45951839145441203   0.281953371838003   0.6778339241356157   0.8408156746392997   0.13184596240883756   0.2682122622912666
0.9972372840383935   0.6467225477192715   0.5581305177390907   0.13596818592323143   0.9706397814650827   0.07192591674001528   0.6375016848789749   0.00852723690202089   0.5767667568905188   0.9987215525024781   0.6971228655573466   0.20521542949326427   0.44531220913659336   0.15601196414300375   0.0776612183163842   0.5604695066117135   0.4201522990832292   0.3248329622368687   0.6181428268619722   0.2785161347737104   0.7423183749476134   0.48401728759756896   0.48629686445313464   0.010303872482443802   0.7450810909092199   0.8372947398782975   0.9281663467140439   0.8743356865592123   0.7744413094441372   0.7653688231382823   0.290664661835069   0.8658084496571915   0.19767455255361838   0.7666472706358042   0.5935417962777224   0.6605930201639272   0.752362343417025   0.6106353064928004   0.5158805779613382   0.1001235135522138   0.3322100443337958   0.2858023442559317   0.897737751099366   0.8216073787785034   0.5898916693861823   0.8017850566583627   0.41144088664623146   0.8113035062960596   0.8448105784769624   0.9644903167800652   0.4832745399321876   0.9369678197368472   0.07036926903282514   0.199121493641783   0.19260987809711858   0.07115937007965574   0.8726947164792067   0.4324742230059789   0.5990680818193961   0.41056634991572855   0.12033237306218172   0.8218389165131784   0.08318750385805784   0.3104428363635147
0.788122328728386   0.5360365722572468   0.18544975275869174   0.48883545758501135   0.19823065934220357   0.734251515598884   0.7740088661124602   0.6775319512889517   0.3534200808652412   0.7697611988188189   0.2907343261802727   0.7405641315521045   0.28305081183241604   0.5706397051770359   0.09812444808315413   0.6694047614724488   0.41035609535320927   0.13816548217105698   0.49905636626375804   0.25883841155672027   0.2900237222910275   0.31632656565787853   0.4158688624057002   0.9483955751932055   0.5019013935626416   0.7802899934006318   0.23041910964700843   0.4595601176081942   0.30367073422043805   0.04603847780174768   0.4564102435345482   0.7820281663192424   0.9502506533551969   0.2762772789829288   0.16567591735427545   0.041464034767137954   0.6671998415227809   0.705637573805893   0.06755146927112134   0.3720592732946892   0.25684374616957156   0.567472091634836   0.5684951030073633   0.11322086173796894   0.966820023878544   0.25114552597695744   0.15262624060166313   0.16482528654476342   0.4649186303159024   0.4708555325763257   0.9222071309546547   0.7052651689365692   0.16124789609546436   0.42481705477457804   0.46579688742010655   0.9232370026173268   0.21099724274026746   0.14853977579164918   0.3001209700658311   0.8817729678501888   0.5437974012174867   0.4429022019857562   0.23256950079470975   0.5097136945554996
0.28695365504791503   0.8754301103509202   0.6640743977873464   0.39649283281753067   0.320133631169371   0.6242845843739627   0.5114481571856833   0.23166754627276726   0.8552150008534686   0.15342905179763708   0.5892410262310286   0.526402377336198   0.6939671047580043   0.7286119970230591   0.12344413881092205   0.6031653747188713   0.4829698620177368   0.5800722212314099   0.8233231687450909   0.7213924068686826   0.9391724608002502   0.13717001924565367   0.5907536679503812   0.21167871231318292   0.6522188057523352   0.2617399088947334   0.9266792701630348   0.8151858794956522   0.33208517458296416   0.6374553245207707   0.41523111297735144   0.583518333222885   0.4768701737294956   0.4840262727231336   0.8259900867463228   0.05711595588668694   0.7829030689714914   0.7554142757000745   0.7025459479354008   0.45395058116781567   0.29993320695375464   0.17534205446866463   0.8792227791903098   0.7325581742991332   0.36076074615350445   0.038172035223010964   0.28846911123992863   0.5208794619859503   0.7085419404011694   0.7764321263282775   0.3617898410768939   0.705693582490298   0.37645676581820514   0.13897680180750685   0.9465587280995424   0.122175249267413   0.8995865920887095   0.6549505290843732   0.12056864135321967   0.06505929338072605   0.11668352311721815   0.8995362533842988   0.4180226934178189   0.6111087122129104
0.8167503161634635   0.7241941989156341   0.5387999142275091   0.8785505379137772   0.45598957000995904   0.6860221636926231   0.2503308029875804   0.35767107592782704   0.7474476296087897   0.9095900373643456   0.8885409619106865   0.6519774934375291   0.3709908637905846   0.7706132355568388   0.9419822338111441   0.5298022441701161   0.4714042717018751   0.11566270647246552   0.8214135924579244   0.46474295078939004   0.35472074858465696   0.21612645308816675   0.4033908990401055   0.8536342385764796   0.5379704324211935   0.4919322541725326   0.8645909848125964   0.9750837006627023   0.08198086241123437   0.8059100904799095   0.614260181825016   0.6174126247348753   0.3345332328024446   0.8963200531155638   0.7257192199143294   0.9654351312973463   0.96354236901186   0.125706817558725   0.7837369861031854   0.4356328871272302   0.49213809730998487   0.01004411108625949   0.962323393645261   0.9708899363378402   0.13741734872532793   0.7939176579980928   0.5589324946051555   0.11725569776136054   0.5994469163041345   0.3019854038255601   0.694341509792559   0.1421719970986582   0.5174660538929001   0.49607531334565064   0.08008132796754307   0.5247593723637829   0.18293282109045553   0.5997552602300869   0.3543621080532136   0.5593242410664366   0.21939045207859553   0.47404844267136187   0.5706251219500282   0.12369135393920647
0.7272523547686106   0.46400433158510235   0.6083017283047673   0.1528014176013663   0.5898350060432828   0.6700866735870097   0.0493692336996117   0.03554571984000576   0.9903880897391483   0.3681012697614495   0.3550277239070526   0.8933737227413475   0.4729220358462481   0.8720259564157988   0.2749463959395096   0.3686143503775647   0.28998921475579253   0.272270696185712   0.920584287886296   0.809290109311128   0.07059876267719702   0.7982222535143502   0.34995916593626775   0.6855987553719216   0.34334640790858634   0.33421792192924776   0.7416574376315006   0.5327973377705553   0.7535114018653036   0.6641312483422381   0.6922882039318888   0.4972516179305495   0.7631233121261555   0.2960299785807886   0.3372604800248362   0.6038778951892019   0.2902012762799073   0.4240040221649898   0.062314084085326654   0.23526354481163725   0.00021206152411477842   0.15173332597927777   0.1417297961990307   0.4259734355005092   0.9296132988469178   0.35351107246492763   0.791770630262763   0.7403746801285876   0.5862668909383314   0.019293150535679884   0.050113192631262356   0.20757734235803238   0.8327554890730278   0.35516190219344174   0.3578249886993735   0.7103257244274829   0.06963217694687232   0.05913192361265313   0.02056450867453727   0.10644782923828093   0.779430900666965   0.6351279014476634   0.9582504245892106   0.8711842844266436
0.7792188391428502   0.4833945754683856   0.8165206283901799   0.4452108489261345   0.8496055402959325   0.12988350300345794   0.024749998127417003   0.7048361687975468   0.26333864935760104   0.11059035246777804   0.9746368054961546   0.49725882643951447   0.43058316028457333   0.7554284502743362   0.6168118167967811   0.7869331020120316   0.360950983337701   0.6962965266616832   0.5962473081222439   0.6804852727737507   0.581520082670736   0.0611686252140198   0.6379968835330333   0.809300988347107   0.8023012435278858   0.5777740497456342   0.8214762551428534   0.3640901394209725   0.9526957032319533   0.44789054674217627   0.7967262570154363   0.6592539706234256   0.6893570538743523   0.3373001942743982   0.8220894515192817   0.16199514418391117   0.258773893589779   0.5818717440000619   0.20527763472250055   0.37506204217187955   0.8978229102520779   0.8855752173383789   0.6090303266002567   0.6945767693981288   0.316302827581342   0.824406592124359   0.9710334430672234   0.8852757810510219   0.5140015840534562   0.24663254237872478   0.14955718792437006   0.5211856416300494   0.5613058808215029   0.7987419956365485   0.3528309309089337   0.8619316710066237   0.8719488269471506   0.46144180136215024   0.530741479389652   0.6999365268227126   0.6131749333573716   0.8795700573620883   0.32546384466715145   0.324874484650833
0.7153520231052937   0.9939948400237095   0.7164335180668948   0.6302977152527042   0.3990491955239516   0.16958824789935048   0.7454000749996714   0.7450219342016823   0.8850476114704954   0.9229557055206257   0.5958428870753013   0.22383629257163284   0.32374173064899253   0.12421370988407722   0.24301195616636764   0.36190462156500913   0.4517929037018419   0.662771908521927   0.7122704767767156   0.6619680947422966   0.8386179703444703   0.7832018511598388   0.3868066321095642   0.33709361009146355   0.12326594723917664   0.7892070111361292   0.6703731140426693   0.7067958948387595   0.724216751715225   0.6196187632367788   0.924973039042998   0.9617739606370772   0.8391691402447297   0.696663057716153   0.32913015196769657   0.7379376680654444   0.5154274095957371   0.5724493478320758   0.08611819580132896   0.3760330465004353   0.06363450589389517   0.9096774393101488   0.37384771902461333   0.7140649517581387   0.22501653554942488   0.1264755881503101   0.9870410869150492   0.3769713416666752   0.10175058831024825   0.3372685770141809   0.3166679728723798   0.6701754468279157   0.37753383659502326   0.7176498137774021   0.39169493382938186   0.7084014861908385   0.5383646963502936   0.02098675606124907   0.06256478186168528   0.9704638181253941   0.022937286754556543   0.44853740822917326   0.9764465860603563   0.5944307716249588
0.9593027808606613   0.5388599689190244   0.602598867035743   0.8803658198668202   0.7342862453112364   0.4123843807687143   0.6155577801206938   0.5033944782001449   0.6325356570009882   0.07511580375453344   0.298889807248314   0.8332190313722293   0.255001820405965   0.35746598997713136   0.9071948734189321   0.1248175451813908   0.7166371240556714   0.33647923391588225   0.8446300915572468   0.15435372705599668   0.6936998373011148   0.887941825686709   0.8681835054968905   0.5599229554310379   0.7343970564404534   0.3490818567676846   0.26558463846114755   0.6795571355642177   0.00011081112921696563   0.9366974759989702   0.6500268583404537   0.17616265736407272   0.3675751541282287   0.8615816722444368   0.3511370510921398   0.3429436259918434   0.11257333372226375   0.5041156822673055   0.44394217767320765   0.21812608081045265   0.3959362096665924   0.16763644835142322   0.5993120861159608   0.06377235375445596   0.7022363723654775   0.2796946226647142   0.7311285806190703   0.5038493983234181   0.9678393159250241   0.9306127658970296   0.4655439421579228   0.8242922627592004   0.9677285047958072   0.9939152898980593   0.815517083817469   0.6481296053951278   0.6001533506675785   0.13233361765362253   0.4643800327253293   0.3051859794032843   0.48758001694531466   0.6282179353863171   0.02043785505212165   0.08705989859283166
0.09164380727872229   0.4605814870348939   0.4211257689361608   0.023287544838375692   0.3894074349132447   0.18088686437017965   0.6899971883170906   0.5194381465149576   0.42156811898822055   0.25027409847315   0.22445324615916779   0.6951458837557571   0.4538396141924134   0.2563588085750907   0.4089361623416987   0.04701627836062938   0.853686263524835   0.12402519092146815   0.9445561296163695   0.7418302989573451   0.3661062465795203   0.4958072555351511   0.9241182745642478   0.6547704003645134   0.274462439300798   0.03522576850025723   0.502992505628087   0.6314828555261377   0.8850550043875532   0.8543389041300776   0.8129953173109964   0.11204470901118017   0.4634868853993327   0.6040648056569276   0.5885420711518287   0.41689882525542304   0.009647271206919321   0.34770599708183686   0.17960590881012992   0.36988254689479366   0.15596100768208435   0.2236808061603687   0.23504977919376047   0.6280522479374486   0.789854761102564   0.7278735506252176   0.31093150462951263   0.9732818475729351   0.5153923218017661   0.6926477821249604   0.8079389990014256   0.3417989920467974   0.6303373174142127   0.8383088779948829   0.9949436816904292   0.22975428303561726   0.16685043201488006   0.23424407233795527   0.4064016105386006   0.8128554577801942   0.15720316080796073   0.8865380752561184   0.2267957017284707   0.44297291088540053
0.0012421531258763846   0.6628572690957497   0.9917459225347103   0.814920662947952   0.2113873920233123   0.9349837184705321   0.6808144179051976   0.8416388153750167   0.6959950702215463   0.24233593634557168   0.872875418903772   0.4998398233282193   0.06565775280733346   0.40402705835068886   0.8779317372133426   0.27008554029260207   0.8988073207924534   0.1697829860127336   0.47153012667474203   0.4572300825124079   0.7416041599844927   0.2832449107566152   0.24473442494627137   0.014257171627007355   0.7403620068586163   0.6203876416608655   0.2529885024115611   0.19933650867905545   0.528974614835304   0.6854039231903334   0.5721740845063635   0.3576976933040387   0.8329795446137577   0.44306798684476173   0.6992986656025916   0.8578578699758194   0.7673217918064242   0.03904092849407286   0.821366928389249   0.5877723296832174   0.8685144710139708   0.8692579424813393   0.3498368017145069   0.13054224717080948   0.1269103110294782   0.5860130317247241   0.10510237676823553   0.11628507554380212   0.3865483041708619   0.9656253900638586   0.8521138743566744   0.9169485668647467   0.857573689335558   0.2802214668735252   0.27993978985031087   0.559250873560708   0.024594144721800226   0.8371534800287636   0.5806411242477193   0.7013930035848885   0.257272352915376   0.7981125515346906   0.7592741958584703   0.11362067390167126
0.38875788190140514   0.9288546090533514   0.4094373941439634   0.9830784267308618   0.26184757087192695   0.3428415773286273   0.3043350173757279   0.8667933511870597   0.8752992667010651   0.37721618726476863   0.4522211430190535   0.949844784322313   0.01772557736550708   0.09699472039124342   0.1722813531687426   0.39059391076160505   0.9931314326437068   0.2598412403624799   0.5916402289210233   0.6892009071767164   0.7358590797283309   0.4617286888277893   0.832366033062553   0.5755802332750451   0.3471011978269258   0.5328740797744379   0.4229286389185896   0.5925018065441834   0.08525362695499883   0.1900325024458106   0.11859362154286172   0.7257084553571237   0.2099543602539338   0.8128163151810419   0.6663724785238082   0.7758636710348107   0.1922287828884267   0.7158215947897986   0.49409112535506566   0.3852697602732057   0.19909735024471986   0.4559803544273186   0.9024508964340423   0.6960688530964892   0.463238270516389   0.9942516655995294   0.07008486337148928   0.12048861982144406   0.11613707268946323   0.4613775858250915   0.6471562244528997   0.5279868132772607   0.0308834457344644   0.27134508337928087   0.528562602910038   0.8022783579201369   0.8209290854805306   0.4585287681982389   0.8621901243862298   0.026414686885326263   0.6287003025921039   0.7427071734084404   0.36809899903116405   0.6411449266121206
0.429602952347384   0.28672681898112173   0.46564810259712175   0.9450760735156314   0.966364681830995   0.2924751533815924   0.39556323922563247   0.8245874536941873   0.8502276091415318   0.831097567556501   0.7484070147727329   0.29660064041692663   0.8193441634070674   0.5597524841772201   0.21984441186269485   0.49432228249678967   0.9984150779265368   0.10122371597898121   0.3576542874764651   0.4679075956114634   0.3697147753344329   0.35851654257054083   0.989555288445301   0.8267626689993428   0.9401118229870489   0.07178972358941908   0.5239071858481793   0.8816865954837114   0.9737471411560539   0.7793145702078267   0.12834394662254678   0.05709914178952416   0.12351953201452208   0.9482170026513257   0.379936931849814   0.7604985013725976   0.3041753686074547   0.3884645184741056   0.16009251998711913   0.2661762188758079   0.30576029068091787   0.2872408024951244   0.8024382325106539   0.7982686232643444   0.936045515346485   0.9287242599245835   0.8128829440653529   0.9715059542650016   0.9959336923594361   0.8569345363351645   0.28897575821717364   0.0898193587812902   0.022186551203382195   0.0776199661273378   0.1606318115946269   0.03272021699176605   0.8986670191888602   0.12940296347601207   0.7806948797448129   0.2722217156191685   0.5944916505814054   0.7409384450019064   0.6206023597576938   0.0060454967433606465
0.28873135990048754   0.4536976425067821   0.8181641272470398   0.2077768734790162   0.35268584455400254   0.5249733825821985   0.005281183181686872   0.23627091921401452   0.35675215219456646   0.668038846247034   0.7163054249645132   0.1464515604327243   0.3345656009911843   0.5904188801196962   0.5556736133698863   0.11373134344095827   0.43589858180232416   0.46101591664368413   0.7749787336250734   0.8415096278217897   0.8414069312209187   0.7200774716417777   0.15437637386737962   0.8354641310784291   0.5526755713204312   0.2663798291349956   0.3362122466203398   0.6276872575994129   0.19998972676642865   0.7414064465527971   0.330931063438653   0.3914163383853984   0.8432375745718621   0.07336760030576307   0.6146256384741398   0.2449647779526741   0.5086719735806778   0.4829487201860668   0.0589520251042534   0.13123343451171582   0.07277339177835368   0.0219328035423827   0.28397329147918   0.2897238066899261   0.23136646055743493   0.30185533190060504   0.12959691761180034   0.45425967561149694   0.6786908892370037   0.03547550276560941   0.7933846709914605   0.826572418012084   0.4787011624705751   0.2940690562128123   0.46245360755280757   0.4351560796266856   0.6354635878987129   0.22070145590704923   0.8478279690786679   0.19019130167401152   0.12679161431803507   0.7377527357209824   0.7888759439744144   0.0589578671622957
0.05401822253968139   0.7158199321785997   0.5049026524952345   0.7692340604723696   0.8226517619822464   0.41396460027799464   0.3753057348834341   0.3149743848608727   0.14396087274524272   0.37848909751238524   0.5819210638919736   0.48840196684878867   0.6652597102746677   0.08442004129957295   0.119467456339166   0.053245887222103036   0.02979612237595472   0.8637185853925238   0.2716394872604982   0.8630545855480916   0.9030045080579197   0.12596584967154134   0.48276354328608373   0.8040967183857958   0.8489862855182383   0.41014591749294166   0.9778608907908493   0.03486265791342619   0.0263345235359918   0.996181317214947   0.6025551559074152   0.7198882730525535   0.882373650790749   0.6176922197025617   0.020634092015441623   0.23148630620376487   0.21711394051608143   0.5332721784029888   0.9011666356762756   0.17824041898166182   0.1873178181401267   0.669553593010465   0.6295271484157775   0.3151858334335703   0.28431331008220706   0.5435877433389237   0.14676360512969372   0.5110891150477744   0.4353270245639688   0.13344182584598208   0.16890271433884443   0.4762264571343483   0.408992501027977   0.1372605086310351   0.5663475584314293   0.7563381840817948   0.5266188502372279   0.5195682889284734   0.5457134664159876   0.5248518778780299   0.3095049097211465   0.9862961105254846   0.644546830739712   0.34661145889636813
0.1221870915810198   0.3167425175150196   0.015019682323934531   0.03142562546279781   0.8378737814988128   0.7731547741760959   0.8682560771942408   0.5203365104150234   0.40254675693484393   0.6397129483301138   0.6993533628553964   0.044110053280675035   0.993554255906867   0.5024524396990787   0.13300580442396714   0.28777186919888026   0.46693540566963904   0.9828841507706053   0.5872923380079795   0.7629199913208503   0.1574304959484925   0.9965880402451207   0.9427455072682676   0.4163085324244822   0.035243404367472725   0.6798455227301011   0.927725824944333   0.38488290696168437   0.19736962286866   0.9066907485540052   0.059469747750092186   0.8645463965466611   0.794822865933816   0.26697780022389145   0.36011638489469583   0.820436343265986   0.8012686100269492   0.7645253605248127   0.22711058047072868   0.5326644740671058   0.33433320435731007   0.7816412097542074   0.6398182424627491   0.7697444827462554   0.17690270840881758   0.7850531695090867   0.6970727351944817   0.3534359503217733   0.14165930404134486   0.10520764677898552   0.7693469102501487   0.9685530433600889   0.9442896811726849   0.19851689822498028   0.7098771625000564   0.1040066468134278   0.14946681523886882   0.9315390980010888   0.3497607776053606   0.2835703035474418   0.3481982052119197   0.16701373747627615   0.12265019713463195   0.750905829480336
0.013865000854609618   0.38537252772206876   0.4828319546718828   0.9811613467340805   0.836962292445792   0.6003193582129821   0.7857592194774011   0.6277253964123073   0.6953029884044472   0.4951117114339966   0.01641230922725256   0.6591723530522184   0.7510133072317623   0.2965948132090164   0.3065351467271961   0.5551657062387907   0.6015464919928936   0.3650557152079275   0.9567743691218356   0.27159540269134885   0.2533482867809738   0.19804197773165136   0.8341241719872036   0.5206895732110128   0.2394832859263642   0.8126694500095826   0.3512922173153208   0.5395282264769323   0.40252099348057213   0.21235009179660044   0.5655329978379195   0.911802830064625   0.707218005076125   0.7172383803626038   0.549120688610667   0.25263047701240654   0.9562046978443626   0.42064356715358747   0.2425855418834709   0.6974647707736159   0.3546582058514691   0.05558785194565996   0.28581117276163537   0.42586936808226705   0.10130991907049529   0.8575458742140086   0.4516870007744318   0.9051797948712542   0.8618266331441311   0.044876424204426016   0.10039478345911106   0.3656515683943219   0.4593056396635589   0.8325263324078256   0.5348617856211915   0.4538487383296969   0.752087634587434   0.11528795204522176   0.9857410970105245   0.20121826131729034   0.7958829367430713   0.6946443848916343   0.7431555551270536   0.5037534905436745
0.44122473089160225   0.6390565329459743   0.4573443823654182   0.0778841224614074   0.339914811821107   0.7815106587319657   0.0056573815909863375   0.17270432759015322   0.4780881786769759   0.7366342345275397   0.9052625981318753   0.8070527591958313   0.01878253901341696   0.9041079021197141   0.3704008125106838   0.35320402086613445   0.266694904425983   0.7888199500744923   0.38465971550015937   0.15198575954884408   0.4708119676829116   0.0941755651828581   0.6415041603731058   0.6482322690051696   0.02958723679130935   0.45511903223688377   0.18415977800768762   0.5703481465437622   0.6896724249702023   0.6736083735049181   0.1785023964167013   0.397643818953609   0.21158424629322647   0.9369741389773784   0.27323979828482603   0.5905910597577777   0.19280170727980953   0.032866236857664176   0.9028389857741422   0.23738703889164325   0.9261068028538265   0.24404628678317178   0.5181792702739829   0.08540127934279917   0.4552948351709149   0.14987072160031367   0.876675109900877   0.43716901033762956   0.4257075983796056   0.6947516893634299   0.6925153318931895   0.8668208637938672   0.7360351734094032   0.02114331585851186   0.5140129354764882   0.4691770448402583   0.5244509271161767   0.08416917688113354   0.24077313719166213   0.8785859850824806   0.3316492198363672   0.051302940023469364   0.3379341514175199   0.6411989461908374
0.4055424169825407   0.8072566532402976   0.819754881143537   0.5557976668480382   0.9502475818116257   0.6573859316399839   0.94307977124266   0.11862865651040863   0.5245399834320201   0.962634242276554   0.25056443934947054   0.25180779271654136   0.788504810022617   0.9414909264180421   0.7365515038729824   0.7826307478762831   0.2640538829064402   0.8573217495369085   0.49577836668132025   0.9040447627938024   0.9324046630700731   0.8060188095134392   0.15784421526380032   0.26284581660296513   0.5268622460875324   0.9987621562731417   0.33808933412026326   0.7070481497549269   0.5766146642759066   0.34137622463315775   0.3950095628776033   0.5884194932445184   0.05207468084388642   0.3787419823566038   0.14444512352813277   0.336611700527977   0.2635698708212694   0.4372510559385616   0.40789361965515036   0.5539809526516939   0.9995159879148292   0.5799293064016531   0.9121152529738301   0.6499361898578915   0.06711132484475618   0.7739104968882138   0.7542710377100298   0.38709037325492635   0.5402490787572238   0.7751483406150722   0.4161817035897666   0.6800422234999994   0.9636344144813173   0.4337721159819144   0.02117214071216329   0.09162273025548111   0.9115597336374308   0.055030133625310645   0.8767270171840306   0.7550110297275041   0.6479898628161613   0.617779077686749   0.46883339752888015   0.2010300770758102
0.6484738749013321   0.037849771285095965   0.55671814455505   0.5510938872179187   0.581362550056576   0.26393927439688214   0.8024471068450202   0.16400351396299234   0.04111347129935216   0.48879093378181   0.3862654032552536   0.4839612904629929   0.07747905681803494   0.05501881779989557   0.3650932625430903   0.39233856020751184   0.16591932318060412   0.999988684174585   0.48836624535905976   0.6373275304800077   0.5179294603644428   0.3822096064878359   0.019532847830179622   0.4362974534041975   0.8694555854631106   0.34435983520273994   0.46281470327512964   0.8852035661862788   0.2880930354065346   0.0804205608058578   0.6603675964301094   0.7212000522232864   0.24697956410718244   0.5916296270240479   0.27410219317485585   0.23723876176029354   0.1695005072891475   0.5366108092241523   0.9090089306317656   0.8449002015527818   0.0035811841085433864   0.5366221250495673   0.42064268527270576   0.20757267107277402   0.48565172374410065   0.1544125185617314   0.40110983744252615   0.7712752176685765   0.6161961382809901   0.8100526833589915   0.9382951341673965   0.8860716514822977   0.3281031028744555   0.7296321225531337   0.27792753773728707   0.16487159925901124   0.08112353876727303   0.13800249552908586   0.0038253445624312245   0.9276328374987177   0.9116230314781255   0.6013916863049336   0.09481641393066567   0.08273263594593597
0.9080418473695822   0.06476956125536629   0.6741737286579599   0.8751599648731619   0.4223901236254815   0.9103570426936348   0.27306389121543373   0.10388474720458542   0.8061939853444915   0.10030435933464339   0.33476875704803716   0.21781309572228771   0.478090882470036   0.37067223678150973   0.056841219310750084   0.05294149646327646   0.39696734370276293   0.23266974125242385   0.053015874748318856   0.12530865896455876   0.4853443122246374   0.6312780549474902   0.9581994608176532   0.04257602301862279   0.5773024648550553   0.566508493692124   0.2840257321596933   0.16741605814546084   0.15491234122957379   0.656151450998489   0.0109618409442596   0.06353131094087543   0.3487183558850823   0.5558470916638457   0.6761930838962225   0.8457182152185877   0.8706274734150463   0.18517485488233598   0.6193518645854723   0.7927767187553113   0.4736601297122834   0.9525051136299121   0.5663359898371535   0.6674680597907525   0.988315817487646   0.3212270586824219   0.6081365290195003   0.6248920367721297   0.4110133526325907   0.754718564990298   0.324110796859807   0.45747597862666883   0.2561010114030169   0.09856711399180884   0.31314895591554737   0.39394466768579345   0.9073826555179345   0.5427200223279631   0.6369558720193249   0.5482264524672057   0.03675518210288819   0.35754516744562714   0.017604007433852605   0.7554497337118945
0.5630950523906048   0.405040053815715   0.4512680175966991   0.08798167392114198   0.5747792349029588   0.08381299513329314   0.8431314885771988   0.4630896371490123   0.16376588227036812   0.3290944301429952   0.5190206917173918   0.005613658522343429   0.9076648708673513   0.23052731615118635   0.20587173580184445   0.61166899083655   0.00028221534941668324   0.6878072938232233   0.5689158637825195   0.0634425383693443   0.9635270332465284   0.33026212637759605   0.5513118563486669   0.3079928046574498   0.40043198085592374   0.925222072561881   0.10004383875196779   0.22001113073630785   0.8256527459529649   0.8414090774285878   0.256912350174769   0.7569214935872955   0.6618868636825967   0.5123146472855927   0.7378916584573771   0.7513078350649521   0.7542219928152456   0.28178733113440635   0.5320199226555327   0.13963884422840214   0.7539397774658289   0.5939800373111831   0.9631040588730132   0.07619630585905786   0.7904127442193004   0.2637179109335871   0.4117922025243463   0.7682035012016081   0.38998076336337667   0.33849583837170605   0.31174836377237847   0.5481923704653001   0.5643280174104117   0.4970867609431182   0.054836013597609506   0.7912708768780046   0.902441153727815   0.9847721136575255   0.3169443551402324   0.039963041813052436   0.14821916091256943   0.7029847825231191   0.7849244324846997   0.9003241975846503
0.3942793834467406   0.10900474521193605   0.8218203736116866   0.8241278917255924   0.6038666392274402   0.8452868342783489   0.4100281710873403   0.055924390523984416   0.21388587586406352   0.5067909959066429   0.0982798073149618   0.5077320200586842   0.6495578584536518   0.009704234963524721   0.0434437937173523   0.7164611431806797   0.7471167047258368   0.024932121305999214   0.72649943857712   0.6764981013676272   0.5988975438132674   0.32194733878288007   0.9415750060924202   0.7761739037829769   0.20461816036652683   0.21294259357094397   0.11975463248073366   0.9520460120573845   0.6007515211390867   0.36765575929259503   0.7097264613933933   0.8961216215334   0.38686564527502315   0.8608647633859521   0.6114466540784316   0.38838960147471585   0.7373077868213713   0.8511605284224274   0.5680028603610793   0.6719284582940361   0.9901910820955345   0.8262284071164282   0.8415034217839593   0.9954303569264089   0.39129353828226715   0.5042810683335481   0.8999284156915391   0.21925645314343203   0.18667537791574035   0.29133847476260416   0.7801737832108055   0.2672104410860475   0.5859238567766537   0.9236827154700091   0.07044732181741212   0.37108881955264744   0.19905821150163056   0.06281795208405702   0.4590006677389805   0.9826992180779316   0.4617504246802592   0.21165742366162965   0.8909978073779012   0.31077075978389546
0.47155934258472465   0.38542901654520145   0.0494943855939419   0.3153404028574865   0.08026580430245746   0.8811479482116533   0.14956596990240273   0.09608394971405447   0.8935904263867172   0.5898094734490492   0.36939218669159724   0.8288735086280069   0.30766656961006345   0.6661267579790401   0.29894486487418515   0.45778468907535946   0.10860835810843288   0.603308805894983   0.8399441971352046   0.47508547099742787   0.6468579334281737   0.3916513822333534   0.9489463897573033   0.1643147112135324   0.17529859084344906   0.006222365688151921   0.8994520041633615   0.8489743083560459   0.09503278654099159   0.12507441747649858   0.7498860342609587   0.7528903586419914   0.2014423601542745   0.5352649440274494   0.38049384756936144   0.9240168500139845   0.8937757905442111   0.8691381860484093   0.08154898269517631   0.466232160938625   0.7851674324357781   0.2658293801534263   0.24160478555997172   0.9911466899411971   0.1383094990076045   0.8741779979200729   0.2926583958026684   0.8268319787276648   0.9630109081641555   0.867955632231921   0.393206391639307   0.9778576703716189   0.8679781216231639   0.7428812147554223   0.6433203573783483   0.22496731172962744   0.6665357614688894   0.207616270727973   0.26282650980898686   0.300950461715643   0.7727599709246783   0.3384780846795637   0.18127752711381054   0.834718300777018
0.9875925384889002   0.07264870452613742   0.9396727415538388   0.8435716108358209   0.8492830394812956   0.19847070660606456   0.6470143457511704   0.016739632108156096   0.8862721313171402   0.33051507437414357   0.25380795411186347   0.03888196173653723   0.018294009693976324   0.5876338596187212   0.6104875967335152   0.8139146500069098   0.35175824822508694   0.3800175888907482   0.3476610869245283   0.5129641882912668   0.5789982773004086   0.04153950421118453   0.16638355981071778   0.6782458875142487   0.5914057388115085   0.9688907996850471   0.22671081825687894   0.834674276678428   0.7421226993302129   0.7704200930789825   0.5796964725057085   0.8179346445702719   0.8558505680130727   0.439905018704839   0.3258885183938451   0.7790526828337346   0.8375565583190964   0.8522711590861177   0.7154009216603299   0.9651380328268249   0.4857983100940094   0.4722535701953695   0.3677398347358016   0.45217384453555803   0.9068000327936008   0.430714065984185   0.20135627492508382   0.7739279570213092   0.3153942939820923   0.4618232662991379   0.9746454566682049   0.9392536803428813   0.5732715946518794   0.6914031732201553   0.39494898416249635   0.12131903577260944   0.7174210266388067   0.2514981545153163   0.06906046576865126   0.3422663529388748   0.8798644683197103   0.3992269954291986   0.35365954410832134   0.37712832011204994
0.39406615822570085   0.9269734252338291   0.9859197093725197   0.9249544755764919   0.4872661254321001   0.49625935924964404   0.7845634344474359   0.15102651855518265   0.17187183145000778   0.03443609295050618   0.8099179777792311   0.21177283821230133   0.5986002367981283   0.3430329197303509   0.4149689936167348   0.0904538024396919   0.8811792101593218   0.09153476521503454   0.3459085278480835   0.7481874495008171   0.0013147418396114437   0.692307769785836   0.9922489837397621   0.3710591293887671   0.6072485836139107   0.7653343445520069   0.006329274367242401   0.4461046538122752   0.11998245818181055   0.26907498530236285   0.22176583991980645   0.29507813525709253   0.9481106267318028   0.23463889235185667   0.41184786214057534   0.08330529704479121   0.3495103899336744   0.8916059726215058   0.9968788685238406   0.9928514946050994   0.4683311797743527   0.8000712074064713   0.6509703406757571   0.24466404510428225   0.46701643793474124   0.1077634376206353   0.658721356935995   0.8736049157155151   0.8597678543208306   0.3424290930686284   0.6523920825687526   0.4275002619032399   0.7397853961390201   0.07335410776626552   0.43062624264894606   0.13242212664614736   0.7916747694072173   0.8387152154144089   0.018778380508370714   0.04911682960135616   0.44216437947354287   0.9471092427929031   0.021899511984530114   0.05626533499625685
0.9738331996991902   0.1470380353864318   0.370929171308773   0.8116012898919747   0.506816761764449   0.0392745977657965   0.7122078143727781   0.9379963741764595   0.6470489074436183   0.6968455046971681   0.05981573180402555   0.5104961122732196   0.9072635113045983   0.6234913969309026   0.6291894891550794   0.3780739856270722   0.11558874189738097   0.7847761815164938   0.6104111086467088   0.328957156025716   0.6734243624238381   0.8376669387235907   0.5885115966621787   0.27269182102945916   0.6995911627246479   0.6906289033371589   0.21758242535340563   0.46109053113748455   0.1927744009601989   0.6513543055713624   0.5053746109806275   0.5230941569610251   0.5457254935165806   0.9545088008741943   0.445558879176602   0.012598044687805527   0.6384619822119824   0.3310174039432917   0.8163693900215225   0.6345240590607333   0.5228732403146014   0.546241222426798   0.20595828137481376   0.3055669030350173   0.8494488778907633   0.7085742837032073   0.6174466847126351   0.03287508200555812   0.14985771516611537   0.017945380366048345   0.3998642593592295   0.5717845508680736   0.9570833142059164   0.36659107479468594   0.894489648378602   0.04869039390704846   0.41135782068933585   0.4120822739204916   0.448930769202   0.03609234921924293   0.7728958384773535   0.08106486997719994   0.6325613791804775   0.4015682901585096
0.2500225981627522   0.534823647550402   0.4266030978056637   0.0960013871234923   0.40057372027198895   0.8262493638471947   0.8091564130930285   0.06312630511793417   0.2507160051058736   0.8083039834811464   0.40929215373379907   0.4913417542498606   0.29363269089995714   0.44171290868646046   0.5148025053551971   0.44265136034281216   0.8822748702106212   0.029630634765968826   0.06587173615319712   0.40655901112356924   0.10937903173326773   0.9485657647887689   0.4333103569727197   0.00499072096505963   0.8593564335705155   0.4137421172383669   0.0067072591670559725   0.9089893338415673   0.4587827132985266   0.5874927533911721   0.1975508460740274   0.8458630287236332   0.208066708192653   0.7791887699100257   0.7882586923402284   0.3545212744737726   0.9144340172926959   0.33747586122356527   0.27345618698503127   0.9118699141309604   0.032159147082074596   0.30784522645759643   0.20758445083183413   0.5053109030073911   0.9227801153488069   0.35927946166882757   0.7742740938591145   0.5003201820423315   0.06342368177829134   0.9455373444304607   0.7675668346920586   0.5913308482007642   0.6046409684797648   0.35804459103928854   0.570015988618031   0.745467819477131   0.39657426028711174   0.5788558211292628   0.7817572962778028   0.39094654500335846   0.4821402429944159   0.24137995990569755   0.5083011092927715   0.4790766308723981
0.4499810959123413   0.9335347334481011   0.30071665846093737   0.9737657278650069   0.5272009805635345   0.5742552717792736   0.5264425646018229   0.4734455458226754   0.4637772987852431   0.6287179273488129   0.7588757299097644   0.8821146976219112   0.8591363303054783   0.27067333630952434   0.1888597412917333   0.1366468781447802   0.4625620700183666   0.6918175151802616   0.40710244501393056   0.7457003331414217   0.9804218270239506   0.45043755527456397   0.8988013357211591   0.2666237022690236   0.5304407311116094   0.5169028218264629   0.5980846772602217   0.2928579744040167   0.0032397505480749327   0.9426475500471893   0.07164211265839883   0.8194124285813413   0.5394624517628318   0.3139296226983764   0.31276638274863444   0.93729773095943   0.6803261214573535   0.04325628638885204   0.12390664145690115   0.8006508528146499   0.21776405143898692   0.3514387712085905   0.7168041964429707   0.05495051967322817   0.23734222441503625   0.9010012159340265   0.8180028607218115   0.7883268174042045   0.7069014933034269   0.38409839410756363   0.21991818346158984   0.49546884300018784   0.703661742755352   0.4414508440603743   0.14827607080319102   0.6760564144188466   0.16419929099252012   0.12752122136199792   0.8355096880545566   0.7387586834594165   0.4838731695351666   0.0842649349731459   0.7116030465976554   0.9381078306447667
0.2661091180961797   0.7328261637645554   0.9947988501546848   0.8831573109715385   0.028766893681143442   0.8318249478305288   0.17679598943287325   0.09483049356733389   0.32186540037771655   0.44772655372296527   0.9568778059712834   0.5993616505671461   0.6182036576223646   0.006275709662590936   0.8086017351680924   0.9233052361482995   0.4540043666298445   0.878754488300593   0.9730920471135358   0.18454655268888298   0.9701311970946779   0.7944895533274471   0.2614890005158804   0.24643872204411635   0.7040220789984982   0.06166338956289172   0.2666901503611956   0.36328141107257794   0.6752551853173547   0.2298384417323628   0.08989416092832235   0.268450917505244   0.3533897849396382   0.7821118880093976   0.13301635495703895   0.669089266938098   0.7351861273172736   0.7758361783468066   0.32441461978894653   0.7457840307897985   0.28118176068742906   0.8970816900462136   0.3513225726754107   0.5612374781009156   0.31105056359275113   0.1025921367187665   0.08983357215953032   0.3147987560567992   0.607028484594253   0.04092874715587478   0.8231434217983347   0.9515173449842212   0.9317732992768981   0.811090305423512   0.7332492608700124   0.6830664274789773   0.57838351433726   0.02897841741411441   0.6002329059129734   0.013977160540879264   0.8431973870199864   0.2531422390673078   0.27581828612402687   0.2681931297510807
0.5620156263325573   0.3560605490210942   0.9244957134486161   0.7069556516501652   0.2509650627398061   0.2534684123023277   0.8346621412890859   0.392156895593366   0.6439365781455532   0.2125396651464529   0.011518719490751122   0.44063955060914467   0.712163278868655   0.40144935972294093   0.27826945862073876   0.7575731231301674   0.13377976453139512   0.37247094230882655   0.6780365527077653   0.7435959625892882   0.29058237751140875   0.11932870324151874   0.40221826658373844   0.4754028328382074   0.7285667511788515   0.7632681542204246   0.4777225531351223   0.7684471811880422   0.4776016884390453   0.5097997419180968   0.6430604118460365   0.3762902855946763   0.8336651102934921   0.29726007677164396   0.6315416923552853   0.9356507349855316   0.12150183142483703   0.8958107170487031   0.3532722337345466   0.17807761185536422   0.9877220668934419   0.5233397747398765   0.6752356810267812   0.4344816492660761   0.6971396893820332   0.4040110714983578   0.2730174144430428   0.9590788164278686   0.9685729382031817   0.6407429172779332   0.7952948613079205   0.19063163523982643   0.4909712497641364   0.13094317535983635   0.15223444946188402   0.8143413496451501   0.6573061394706443   0.8336830985881923   0.5206927571065987   0.8786906146596185   0.5358043080458073   0.9378723815394893   0.1674205233720521   0.7006130028042543
0.5480822411523654   0.4145326067996128   0.4921848423452709   0.2661313535381782   0.8509425517703322   0.010521535301255026   0.21916742790222807   0.30705253711030955   0.8823696135671505   0.3697786180233218   0.42387256659430755   0.11642090187048311   0.39139836380301407   0.23883544266348547   0.27163811713242353   0.302079552225333   0.7340922243323698   0.4051523440752931   0.7509453600258248   0.4233889375657145   0.1982879162865625   0.4672799625358038   0.5835248366537727   0.7227759347614602   0.6502056751341971   0.05274735573619099   0.09133999430850187   0.456644581223282   0.799263123363865   0.042225820434935966   0.8721725664062738   0.14959204411297244   0.9168935097967145   0.6724472024116142   0.4482999998119663   0.03317114224248933   0.5254951459937003   0.4336117597481287   0.17666188267954275   0.7310915900171564   0.7914029216613305   0.028459415672835574   0.4257165226537179   0.30770265245144185   0.593115005374768   0.5611794531370318   0.8421916859999452   0.5849267176899817   0.9429093302405709   0.5084320974008408   0.7508516916914433   0.1282821364666997   0.143646206876706   0.46620627696590483   0.8786791252851694   0.9786900923537273   0.2267526970799916   0.7937590745542906   0.43037912547320323   0.9455189501112379   0.7012575510862913   0.36014731480616197   0.2537172427936605   0.21442736009408156
0.9098546294249606   0.3316878991333264   0.8280007201399426   0.9067247076426397   0.3167396240501926   0.7705084459962946   0.9858090341399974   0.321797989952658   0.3738302938096217   0.2620763485954538   0.2349573424485541   0.19351585348595832   0.23018408693291567   0.795870071629549   0.3562782171633846   0.2148257611322311   0.0034313898529240725   0.0021109970752583467   0.9258990916901814   0.2693068110209932   0.30217383876663284   0.6419636822690964   0.6721818488965209   0.054879450926911606   0.39231920934167214   0.31027578313577   0.8441811287565782   0.14815474328427192   0.07557958529147953   0.5397673371394753   0.8583720946165809   0.8263567533316138   0.7017492914818578   0.2776909885440215   0.6234147521680268   0.6328408998456555   0.4715652045489422   0.4818209169144725   0.2671365350046422   0.4180151387134245   0.4681338146960181   0.4797099198392141   0.3412374433144608   0.1487083276924313   0.1659599759293853   0.8377462375701178   0.6690555944179399   0.0938288767655197   0.7736407665877132   0.5274704544343478   0.8248744656613616   0.9456741334812477   0.6980611812962336   0.9877031172948725   0.9665023710447808   0.1193173801496339   0.9963118898143758   0.710012128750851   0.34308761887675393   0.48647648030397833   0.5247466852654336   0.22819121183637847   0.07595108387211175   0.06846134159055388
0.056612870569415455   0.7484812919971643   0.734713640557651   0.9197530138981226   0.8906528946400302   0.9107350544270465   0.06565804613971103   0.8259241371326029   0.117012128052317   0.38326459999269874   0.24078358047834944   0.8802500036513551   0.4189509467560834   0.39556148269782626   0.2742812094335687   0.7609326235017212   0.4226390569417076   0.6855493539469752   0.9311935905568148   0.27445614319774286   0.897892371676274   0.45735814211059683   0.855242506684703   0.205994801607189   0.8412795011068586   0.7088768501134325   0.12052886612705212   0.2862417877090664   0.9506266064668284   0.798141795686386   0.05487081998734108   0.4603176505764635   0.8336144784145114   0.41487719569368725   0.8140872395089916   0.5800676469251084   0.414663531658428   0.019315712995860986   0.5398060300754229   0.8191350234233872   0.9920244747167204   0.3337663590488857   0.6086124395186081   0.5446788802256444   0.09413210304044639   0.8764082169382889   0.7533699328339051   0.33868407861845534   0.25285260193358783   0.1675313668248564   0.6328410667068529   0.05244229090938895   0.3022259954667594   0.36938957113847043   0.5779702467195119   0.5921246403329254   0.468611517052248   0.9545123754447832   0.7638830072105203   0.012056993407817004   0.05394798539381997   0.9351966624489222   0.2240769771350973   0.1929219699844298
0.06192351067709955   0.6014303034000366   0.6154645376164892   0.6482430897587854   0.9677914076366532   0.7250220864617476   0.8620946047825842   0.3095590111403301   0.7149388057030653   0.5574907196368912   0.22925353807573112   0.2571167202309411   0.41271281023630596   0.1881011484984208   0.6512832913562192   0.6649920798980157   0.944101293184058   0.2335887730536376   0.887400284145699   0.6529350864901987   0.890153307790238   0.2983921106047154   0.6633233070106017   0.4600131165057689   0.8282297971131385   0.6969618072046788   0.04785876939411253   0.8117700267469835   0.8604383894764853   0.9719397207429312   0.18576416461152842   0.5022110156066534   0.14549958377341993   0.41444900110604   0.9565106265357973   0.24509429537571226   0.732786773537114   0.2263478526076192   0.30522733517957806   0.5801022154776966   0.788685480353056   0.9927590795539816   0.417827051033879   0.9271671289874979   0.898532172562818   0.6943669689492662   0.7545037440232774   0.467154012481729   0.07030237544967957   0.9974051617445874   0.7066449746291648   0.6553839857347455   0.20986398597319428   0.025465441001656142   0.5208808100176364   0.1531729701280921   0.06436440219977435   0.6110164398956162   0.5643701834818391   0.9080786747523798   0.3315776286626604   0.38466858728799697   0.25914284830226103   0.3279764592746833
0.5428921483096043   0.39190950773401534   0.841315797268382   0.4008093302871854   0.6443599757467863   0.6975425387847491   0.08681205324510466   0.9336553178054564   0.5740576002971067   0.7001373770401618   0.38016707861593985   0.2782713320707109   0.36419361432391245   0.6746719360385056   0.8592862685983035   0.12509836194261878   0.2998292121241381   0.06365549614288944   0.29491608511646444   0.21701968719023892   0.9682515834614778   0.6789869088548925   0.03577323681420339   0.8890432279155557   0.4253594351518734   0.28707740112087715   0.1944574395458214   0.4882338976283703   0.7809994594050871   0.5895348623361281   0.10764538630071674   0.5545785798229138   0.20694185910798035   0.8893974852959663   0.7274783076847768   0.27630724775220294   0.8427482447840678   0.21472554925746073   0.8681920390864734   0.15120888580958414   0.5429190326599298   0.15107005311457128   0.573275953970009   0.9341891986193452   0.574667449198452   0.4720831442596788   0.5375027171558056   0.04514597070378955   0.14930801404657865   0.18500574313880164   0.3430452776099842   0.5569120730754192   0.3683085546414916   0.5954708808026736   0.23539989130926744   0.0023334932525054444   0.16136669553351124   0.7060733955067072   0.5079215836244906   0.7260262455003025   0.31861845074944334   0.4913478462492465   0.6397295445380172   0.5748173596907183
0.7756994180895136   0.3402777931346752   0.0664535905680082   0.6406281610713732   0.2010319688910615   0.8681946488749964   0.5289508734122026   0.5954821903675837   0.05172395484448286   0.6831889057361948   0.18590559580221844   0.038570117292164335   0.6834154002029913   0.08771802493352122   0.950505704492951   0.036236624039658896   0.5220487046694801   0.381644629426814   0.44258412086846044   0.3102103785393564   0.20343025392003672   0.8902967831775674   0.8028545763304432   0.7353930188486381   0.4277308358305231   0.5500189900428922   0.7364009857624351   0.09476485777726484   0.22669886693946165   0.6818243411678958   0.20745011235023242   0.49928266740968125   0.17497491209497879   0.998635435431701   0.021544516548013988   0.4607125501175169   0.4915595118919875   0.9109174104981798   0.071038812055063   0.424475926077858   0.9695108072225074   0.5292727810713658   0.6284546911866026   0.11426554753850161   0.7660805533024707   0.6389759978937983   0.8256001148561594   0.3788725286898636   0.3383497174719476   0.08895700785090609   0.08919912909372428   0.28410767091259875   0.11165085053248593   0.4071326666830103   0.8817490167434918   0.7848250035029175   0.9366759384375072   0.40849723125130927   0.8602045001954779   0.3241124533854007   0.4451164265455197   0.4975798207531295   0.7891656881404149   0.8996365273075426
0.47560561932301226   0.9683070396817637   0.1607109969538123   0.785370979769041   0.7095250660205416   0.3293310417879654   0.335110882097653   0.4064984510791774   0.37117534854859396   0.24037403393705933   0.2459117530039287   0.12239078016657869   0.25952449801610805   0.8332413672540491   0.3641627362604368   0.33756577666366117   0.3228485595786009   0.42474413600273975   0.5039582360649589   0.013453323278260498   0.8777321330330813   0.9271643152496102   0.714792547924544   0.11381679597071784   0.40212651371006897   0.9588572755678465   0.5540815509707318   0.3284458162016768   0.6926014476895275   0.629526233779881   0.2189706688730788   0.9219473651224993   0.3214260991409335   0.38915219984282173   0.9730589158691502   0.7995565849559206   0.061901601124825435   0.5559108325887727   0.6088961796087133   0.46199080829225947   0.7390530415462245   0.13116669658603297   0.10493794354375433   0.448537485013999   0.8613209085131432   0.20400238133642273   0.39014539561921024   0.33472068904328117   0.4591943948030743   0.24514510576857626   0.8360638446484785   0.006274872841604374   0.7665929471135469   0.6156188719886951   0.6170931757753997   0.08432750771910504   0.44516684797261336   0.22646667214587343   0.6440342599062495   0.2847709227631844   0.3832652468477879   0.6705558395571007   0.035138080297536255   0.8227801144709249
0.6442122053015634   0.5393891429710678   0.9302001367537819   0.37424262945692593   0.7828912967884201   0.335386761634645   0.5400547411345716   0.03952194041364476   0.3236969019853458   0.09024165586606872   0.7039908964860933   0.033247067572040385   0.557103954871799   0.47462278387737356   0.08689772071069356   0.9489195598529353   0.1119371068991856   0.24815611173150012   0.442863460804444   0.6641486370897509   0.7286718600513977   0.5776002721743995   0.40772538050690776   0.841368522618826   0.08445965474983427   0.0382111292033317   0.4775252437531258   0.4671258931619001   0.3015683579614142   0.7028243675686867   0.9374705026185541   0.42760395274825536   0.9778714559760684   0.612582711702618   0.23347960613246094   0.394356885176215   0.4207675011042694   0.13795992782524444   0.1465818854217674   0.4454373253232796   0.30883039420508385   0.8898038160937444   0.7037184246173234   0.7812886882335287   0.5801585341536861   0.3122035439193449   0.2959930441104156   0.9399201656147026   0.4956988794038519   0.2739924147160132   0.8184678003572898   0.47279427245280253   0.1941305214424377   0.5711680471473265   0.8809972977387356   0.04519031970454717   0.21625906546636933   0.9585853354447085   0.6475176916062747   0.6508334345283322   0.7954915643620999   0.820625407619464   0.5009358061845073   0.20539610920505258
0.4866611701570161   0.9308215915257196   0.7972173815671839   0.4241074209715239   0.9065026360033299   0.6186180476063748   0.5012243374567683   0.4841872553568213   0.41080375659947804   0.34462563289036163   0.6827565370994785   0.01139298290401873   0.21667323515704037   0.7734575857430351   0.8017592393607429   0.9662026631994716   0.0004141696906710345   0.8148722502983267   0.15424154775446822   0.31536922867113937   0.20492260532857112   0.9942468426788627   0.6533057415699609   0.10997311946608677   0.718261435171555   0.06342525115314299   0.856088360002777   0.6858656984945629   0.8117587991682251   0.44480720354676817   0.3548640225460087   0.2016784431377416   0.40095504256874703   0.10018157065640657   0.6721074854465302   0.1902854602337229   0.18428180741170666   0.3267239849133714   0.8703482460857873   0.22408279703425132   0.18386763772103562   0.5118517346150447   0.716106698331319   0.908713568363112   0.9789450323924646   0.5176048919361821   0.06280095676135813   0.7987404488970252   0.26068359722090945   0.4541796407830391   0.20671259675858114   0.11287475040246231   0.44892479805268437   0.00937243723627086   0.8518485742125724   0.9111963072647207   0.047969755483937365   0.9091908665798643   0.17974108876604228   0.7209108470309978   0.8636879480722307   0.5824668816664929   0.30939284268025496   0.49682804999674646
0.6798203103511951   0.07061514705144815   0.5932861443489359   0.5881144816336344   0.7008752779587306   0.5530102551152661   0.5304851875875778   0.7893740327366093   0.4401916807378211   0.09883061433222706   0.3237725908289967   0.676499282334147   0.9912668826851367   0.0894581770959562   0.47192401661642425   0.7653029750694263   0.9432971272011994   0.1802673105160919   0.29218292785038197   0.044392128038428506   0.07960917912896867   0.597800428849599   0.982790085170127   0.5475640780416821   0.3997888687777736   0.5271852817981509   0.38950394082119105   0.9594495964080475   0.698913590819043   0.9741750266828848   0.8590187532336132   0.17007556367143822   0.25872191008122186   0.8753444123506577   0.5352461624046165   0.49357628133729126   0.2674550273960851   0.7858862352547015   0.06332214578819235   0.7282733062678649   0.3241579001948858   0.6056189247386096   0.7711392179378104   0.6838811782294364   0.2445487210659171   0.007818495889010565   0.7883491327676835   0.1363171001877544   0.8447598522881435   0.4806332140908597   0.39884519194649243   0.17686750377970684   0.1458462614691005   0.5064581874079749   0.5398264387128792   0.006791940108268615   0.8871243513878786   0.6311137750573171   0.004580276308262583   0.5132156587709774   0.6196693239917935   0.8452275398026157   0.9412581305200702   0.7849423525031124
0.29551142379690776   0.23960861506400602   0.1701189125822598   0.10106117427367602   0.05096270273099064   0.23179011917499545   0.3817697798145764   0.9647440740859217   0.20620285044284714   0.7511569050841358   0.982924587868084   0.7878765703062148   0.060356588973746614   0.24469871767616092   0.4430981491552048   0.7810846301979462   0.17323223758586798   0.6135849426188438   0.4385178728469422   0.2678689714269688   0.5535629135940745   0.7683574028162281   0.49725974232687203   0.48292661892385635   0.25805148979716674   0.5287487877522221   0.32714082974461217   0.3818654446501803   0.2070887870661761   0.29695866857722664   0.9453710499300358   0.4171213705642587   0.0008859366233289528   0.5458017634930908   0.9624464620619518   0.6292448002580439   0.9405293476495823   0.3011030458169299   0.519348312906747   0.8481601700600977   0.7672971100637144   0.6875181031980862   0.08083044005980478   0.580291198633129   0.2137341964696399   0.919160700381858   0.5835706977329328   0.09736457970927259   0.9556827066724731   0.390411912629636   0.25642986798832057   0.7154991350590922   0.7485939196062971   0.09345324405240935   0.3110588180582848   0.2983777644948336   0.7477079829829681   0.5476514805593184   0.34861235599633295   0.6691329642367897   0.8071786353333859   0.24654843474238858   0.8292640430895859   0.8209727941766919
0.03988152526967143   0.5590303315443024   0.7484336030297811   0.240681595543563   0.8261473288000315   0.6398696311624443   0.16486290529684838   0.1433170158342904   0.8704646221275584   0.24945771853280835   0.9084330373085278   0.4278178807751981   0.12187070252126125   0.156004474480399   0.597374219250243   0.12944011628036456   0.3741627195382931   0.6083529939210806   0.24876186325391006   0.46030715204357486   0.5669840842049073   0.3618045591786919   0.41949782016432413   0.639334357866883   0.5271025589352358   0.8027742276343895   0.671064217134543   0.3986527623233199   0.7009552301352043   0.16290459647194525   0.5062013118376946   0.2553357464890295   0.830490608007646   0.9134468779391369   0.5977682745291668   0.8275178657138313   0.7086199054863848   0.7574424034587379   0.0003940552789237525   0.6980777494334668   0.33445718594809165   0.14908940953765737   0.7516321920250137   0.23777059738989195   0.7674731017431844   0.7872848503589654   0.33213437186068956   0.5984362395230091   0.24037054280794848   0.9845106227245759   0.6610701547261466   0.1997834771996891   0.5394153126727441   0.8216060262526307   0.15486884288845207   0.9444477307106596   0.7089247046650982   0.9081591483134938   0.5571005683592853   0.1169298649968282   0.0003047991787133537   0.15071674485475586   0.5567065130803616   0.4188521155633614
0.6658476132306217   0.0016273353170985017   0.8050743210553478   0.1810815181734694   0.8983745114874374   0.21434248495813307   0.47293994919465826   0.5826452786504603   0.6580039686794888   0.22983186223355723   0.8118697944685116   0.38286180145077126   0.11858865600674477   0.4082258359809266   0.6570009515800596   0.4384140707401117   0.4096639513416467   0.5000666876674329   0.09990038322077428   0.32148420574328346   0.40935915216293334   0.34934994281267695   0.5431938701404128   0.9026320901799221   0.7435115389323116   0.3477226074955785   0.7381195490850649   0.7215505720064527   0.8451370274448743   0.13338012253744538   0.2651795998904066   0.13890529335599233   0.18713305876538536   0.9035482603038881   0.453309805421895   0.756043491905221   0.06854440275864057   0.4953224243229616   0.7963088538418354   0.3176294211651094   0.6588804514169939   0.9952557366555288   0.6964084706210611   0.996145215421826   0.2495212992540606   0.6459057938428517   0.1532146004806484   0.09351312524190387   0.506009760321749   0.2981831863472733   0.4150950513955835   0.3719625532354512   0.6608727328768748   0.1648030638098279   0.14991545150517688   0.23305725987945886   0.4737396741114894   0.2612548035059397   0.6966056460832819   0.4770137679742378   0.40519527135284883   0.7659323791829782   0.9002967922414464   0.15938434680912836
0.7463148199358549   0.7706766425274494   0.20388832162038534   0.1632391313873024   0.4967935206817943   0.1247708486845976   0.050673721139736956   0.06972600614539853   0.9907837603600453   0.8265876623373243   0.6355786697441534   0.6977634529099473   0.3299110274831706   0.6617845985274964   0.4856632182389766   0.4647061930304885   0.8561713533716812   0.40052979502155667   0.7890575721556947   0.9876924250562507   0.4509760820188324   0.6345974158385785   0.8887607799142483   0.8283080782471224   0.7046612620829774   0.8639207733111292   0.6848724582938629   0.6650689468598199   0.20786774140118316   0.7391499246265315   0.634198737154126   0.5953429407144214   0.21708398104113785   0.9125622622892072   0.9986200674099724   0.897579487804474   0.8871729535579673   0.25077766376171085   0.5129568491709959   0.43287329477398556   0.03100160018628612   0.8502478687401541   0.7238992770153012   0.44518086971773485   0.5800255181674537   0.21565045290157564   0.8351384971010529   0.6168727914706126   0.8753642560844763   0.3517296795904465   0.15026603880719   0.9518038446107926   0.6674965146832932   0.6125797549639149   0.516067301653064   0.35646090389637125   0.4504125336421553   0.7000174926747077   0.5174472342430916   0.4588814160918972   0.563239580084188   0.4492398289129969   0.004490385072095659   0.02600812131791163
0.5322379798979019   0.5989919601728427   0.2805911080567945   0.5808272516001768   0.9522124617304482   0.3833415072712671   0.44545261095574157   0.9639544601295642   0.0768482056459718   0.031611827680820624   0.29518657214855154   0.012150615518771606   0.40935169096267865   0.4190320727169057   0.7791192704954875   0.6556897116224004   0.9589391573205234   0.719014580042198   0.26167203625239593   0.1968082955305032   0.3956995772363354   0.2697747511292011   0.2571816511803003   0.17080017421259155   0.8634615973384335   0.6707827909563583   0.9765905431235058   0.5899729226124147   0.9112491356079854   0.2874412836850912   0.5311379321677643   0.6260184624828505   0.8344009299620136   0.2558294560042706   0.23595136001921269   0.6138678469640789   0.42504923899933494   0.8367973832873649   0.4568320895237252   0.9581781353416786   0.4661100816788115   0.11778280324516696   0.1951600532713293   0.7613698398111755   0.07041050444247614   0.8480080521159659   0.937978402091029   0.5905696655985838   0.2069489071040426   0.17722526115960757   0.9613878589675232   0.0005967429861690506   0.2956997714960572   0.8897839774745163   0.430249926799759   0.3745782805033185   0.46129884153404355   0.6339545214702458   0.1942985667805463   0.7607104335392395   0.03624960253470864   0.7971571381828809   0.7374664772568211   0.8025322981975609
0.5701395208558971   0.6793743349377139   0.5423064239854918   0.04116245838638553   0.49972901641342093   0.8313662828217481   0.6043280218944628   0.4505927927878017   0.29278010930937837   0.6541410216621404   0.6429401629269396   0.4499960498016326   0.9970803378133212   0.7643570441876241   0.21269023612718058   0.07541776929831415   0.5357814962792776   0.1304025227173783   0.018391669346634294   0.3147073357590746   0.49953189374456897   0.3332453845344974   0.2809251920898132   0.5121750375615137   0.9293923728886719   0.6538710495967835   0.7386187681043214   0.4710125791751282   0.42966335647525095   0.8225047667750355   0.13429074620985862   0.0204197863873265   0.13688324716587255   0.16836374511289506   0.49135058328291903   0.5704237365856939   0.13980290935255138   0.40400670092527097   0.27866034715573845   0.4950059672873797   0.6040214130732737   0.2736041782078927   0.2602686778091042   0.1802986315283051   0.10448951932870477   0.9403587936733953   0.979343485719291   0.6681235939667914   0.17509714644003288   0.2864877440766117   0.24072471761496955   0.1971110147916632   0.7454337899647819   0.4639829773015762   0.10643397140511093   0.1766912284043367   0.6085505427989094   0.2956192321886812   0.6150833881221919   0.6062674918186428   0.468747633446358   0.8916125312634102   0.3364230409664535   0.11126152453126312
0.8647262203730842   0.6180083530555175   0.0761543631573493   0.930962893002958   0.7602367010443795   0.6776495593821222   0.09681087743805836   0.2628392990361666   0.5851395546043466   0.39116181530551053   0.8560861598230888   0.0657282842445034   0.8397057646395646   0.9271788380039343   0.7496521884179779   0.8890370558401667   0.23115522184065523   0.6315596058152532   0.13456880029578597   0.28276956402152387   0.7624075883942972   0.7399470745518429   0.7981457593293325   0.17150803949026072   0.8976813680212129   0.12193872149632545   0.7219913961719832   0.2405451464873027   0.13744466697683344   0.4442891621142032   0.6251805187339249   0.9777058474511361   0.5523051123724868   0.05312734680869268   0.769094358910836   0.9119775632066327   0.7125993477329222   0.12594850880475839   0.019442170492858166   0.022940507366465992   0.481444125892267   0.4943889029895053   0.8848733701970722   0.7401709433449422   0.7190365374979698   0.7544418284376623   0.08672761086773968   0.5686629038546814   0.8213551694767569   0.6325031069413368   0.36473621469575646   0.3281177573673787   0.6839105024999235   0.18821394482713366   0.7395556959618316   0.3504119099162426   0.13160539012743658   0.135086598018441   0.9704613370509956   0.43843434670960996   0.41900604239451433   0.009138089213682603   0.9510191665581375   0.41549383934314393
0.9375619165022473   0.5147491862241773   0.06614579636106521   0.6753228959982018   0.21852537900427754   0.760307357786515   0.9794181854933255   0.10665999214352039   0.39717020952752063   0.12780425084517816   0.614681970797569   0.7785422347761417   0.7132597070275972   0.9395903060180445   0.8751262748357375   0.42813032485989905   0.5816543169001607   0.8045037079996035   0.9046649377847419   0.9896959781502891   0.16264827450564628   0.7953656187859209   0.9536457712266044   0.5742021388071451   0.22508635800339893   0.28061643256174357   0.8874999748655392   0.8988792428089434   0.006560978999121397   0.5203090747752286   0.9080817893722137   0.792219250665423   0.6093907694716008   0.3925048239300504   0.29339981857464464   0.0136770158892813   0.8961310624440035   0.4529145179120059   0.4182735437389072   0.5855466910293823   0.31447674554384286   0.6484108099124024   0.5136086059541654   0.5958507128790932   0.1518284710381966   0.8530451911264815   0.5599628347275608   0.02164857407194799   0.9267421130347977   0.5724287585647378   0.6724628598620216   0.12276933126300464   0.9201811340356763   0.052119683789509354   0.7643810704898079   0.3305500805975817   0.31079036456407555   0.659614859859459   0.47098125191516327   0.31687306470830034   0.414659302120072   0.20670034194745313   0.05270770817625606   0.7313263736789181
0.10018255657622913   0.5582895320350507   0.5390991022220908   0.13547566079982495   0.9483540855380326   0.7052443409085694   0.9791362674945299   0.11382708672787697   0.021611972503234874   0.13281558234383142   0.3066734076325083   0.9910577554648723   0.10143083846755861   0.08069589855432206   0.5422923371427004   0.6605076748672907   0.7906404739034831   0.4210810386948631   0.07131108522753712   0.34363461015899033   0.37598117178341106   0.21438069674740995   0.01860337705128106   0.6123082364800722   0.27579861520718196   0.6560911647123592   0.47950427482919034   0.47683257568024723   0.32744452966914944   0.9508468238037899   0.5003680073346605   0.3630054889523702   0.30583255716591456   0.8180312414599584   0.19369459970215216   0.37194773348749793   0.20440171869835594   0.7373353429056364   0.6514022625594518   0.7114400586202072   0.41376124479487286   0.31625430421077333   0.5800911773319147   0.36780544846121693   0.03778007301146176   0.10187360746336335   0.5614878002806336   0.7554972119811447   0.7619814578042798   0.44578244275100415   0.0819835254514433   0.2786646363008975   0.4345369281351304   0.4949356189472143   0.5816155181167828   0.9156591473485273   0.12870437096921583   0.6769043774872558   0.38792091841463067   0.5437114138610294   0.92430265227086   0.9395690345816194   0.7365186558551788   0.8322713552408221
0.5105414074759871   0.6233147303708462   0.1564274785232642   0.4644659067796052   0.4727613344645253   0.5214411229074828   0.5949396782426305   0.7089686947984605   0.7107798766602454   0.07565868015647861   0.5129561527911872   0.4303040584975629   0.2762429485251151   0.5807230612092643   0.9313406346744044   0.5146449111490357   0.14753857755589928   0.9038186837220085   0.5434197162597737   0.9709334972880064   0.22323592528503938   0.964249649140389   0.8069010604045949   0.13866214204718424   0.7126945178090524   0.3409349187695429   0.6504735818813306   0.6741962352675791   0.239933183344527   0.8194937958620602   0.0555339036387001   0.9652275404691186   0.5291533066842815   0.7438351157055815   0.5425777508475128   0.5349234819715557   0.2529103581591664   0.16311205449631716   0.6112371161731085   0.02027857082251996   0.10537178060326716   0.2592933707743087   0.06781739991333476   0.04934507353451362   0.8821358553182278   0.2950437216339196   0.26091633950873994   0.9106829314873294   0.16944133750917545   0.9541088028643767   0.6104427576274093   0.23648669621975033   0.9295081541646485   0.1346150070023166   0.5549088539887091   0.27125915575063175   0.4003548474803669   0.39077989129673507   0.012331103141196304   0.736335673779076   0.14744448932120047   0.2276678368004179   0.40109398696808785   0.7160571029565561
0.04207270871793332   0.9683744660261092   0.3332765870547531   0.6667120294220426   0.15993685339970554   0.6733307443921897   0.07236024754601318   0.7560290979347131   0.9904955158905301   0.7192219415278129   0.46191748991860393   0.5195424017149628   0.060987361725881636   0.5846069345254963   0.9070086359298948   0.24828324596433105   0.6606325142455147   0.1938270432287612   0.8946775327886984   0.511947572185255   0.5131880249243143   0.9661592064283433   0.49358354582061065   0.7958904692286989   0.4711153162063809   0.9977847404022341   0.16030695876585752   0.12917843980665636   0.3111784628066754   0.32445399601004443   0.08794671121984435   0.3731493418719432   0.3206829469161453   0.6052320544822315   0.6260292213012404   0.8536069401569805   0.2596955851902637   0.020625119956735227   0.7190205853713456   0.6053236941926494   0.599063070944749   0.826798076727974   0.8243430525826472   0.0933761220073944   0.08587504602043469   0.8606388702996307   0.3307595067620365   0.29748565277869554   0.6147597298140538   0.8628541298973967   0.170452547996179   0.16830721297203918   0.30358126700737836   0.5384001338873523   0.08250583677633468   0.795157871100096   0.982898320091233   0.9331680794051208   0.45647661547509427   0.9415509309431155   0.7232027349009693   0.9125429594483856   0.7374560301037486   0.3362272367504661
0.12413966395622039   0.08574488272041153   0.9131129775211014   0.24285111474307175   0.03826461793578571   0.2251060124207808   0.5823534707590649   0.9453654619643762   0.4235048881217319   0.3622518825233841   0.41190092276288587   0.777058248992337   0.11992362111435359   0.8238517486360317   0.3293950859865512   0.981900377892241   0.13702530102312055   0.890683669230911   0.8729184705114569   0.040349446949125525   0.4138225661221512   0.9781407097825254   0.1354624404077083   0.7041222101986594   0.2896829021659308   0.8923958270621138   0.22234946288660687   0.46127109545558764   0.2514182842301451   0.6672898146413331   0.639995992127542   0.5159056334912114   0.8279133961084132   0.30503793211794905   0.2280950693646561   0.7388473844988744   0.7079897749940596   0.4811861834819173   0.8986999833781049   0.7569470066066334   0.570964473970939   0.5905025142510063   0.025781512866647975   0.7165975596575078   0.15714190784878782   0.6123618044684809   0.8903190724589397   0.012475349458848477   0.867459005682857   0.719965977406367   0.6679696095723329   0.5512042540032609   0.6160407214527119   0.052676162765033875   0.027973617444790856   0.03529862051204941   0.7881273253442987   0.7476382306470848   0.7998785480801348   0.29645123601317497   0.0801375503502392   0.26645204716516757   0.9011785647020298   0.5395042294065416
0.5091730763793002   0.6759495329141613   0.8753970518353819   0.8229066697490337   0.35203116853051236   0.06358772844568039   0.9850779793764423   0.8104313202901853   0.48457216284765536   0.3436217510393134   0.3171083698041094   0.25922706628692443   0.8685314413949434   0.2909455882742795   0.28913475235931857   0.22392844577487503   0.0804041160506447   0.5433073576271947   0.48925620427918376   0.9274772097617   0.0002665657004055004   0.27685531046202716   0.5880776395771539   0.3879729803551584   0.4910934893211053   0.6009057775478659   0.712680587741772   0.5650663106061247   0.13906232079059294   0.5373180491021855   0.7276026083653299   0.7546349903159394   0.6544901579429376   0.19369629806287209   0.4104942385612204   0.49540792402901496   0.7859587165479941   0.9027507097885925   0.12135948620190186   0.2714794782541399   0.7055546004973494   0.35944335216139783   0.632103281922718   0.3440022684924399   0.7052880347969439   0.08258804169937073   0.04402564234556416   0.9560292881372815   0.2141945454758386   0.48168226415150484   0.33134505460379216   0.39096297753115683   0.07513222468524566   0.9443642150493193   0.6037424462384623   0.6363279872152174   0.4206420667423081   0.7506679169864473   0.1932482076772419   0.14092006318620248   0.634683350194314   0.8479172071978547   0.07188872147534005   0.8694405849320626
0.9291287496969646   0.48847385503645685   0.43978543955262195   0.5254383164396227   0.22384071490002058   0.4058858133370862   0.3957597972070578   0.5694090283023412   0.009646169424181972   0.9242035491855813   0.06441474260326568   0.17844605077118433   0.9345139447389363   0.9798393341362619   0.46067229636480334   0.5421180635559669   0.5138718779966283   0.22917141714981465   0.26742408868756146   0.40119800036976444   0.8791885278023143   0.3812542099519599   0.1955353672122214   0.5317574154377019   0.9500597781053497   0.892780354915503   0.7557499276595995   0.006319098998079279   0.7262190632053291   0.4868945415784169   0.35999013045254163   0.4369100706957381   0.7165728937811472   0.5626909923928356   0.29557538784927595   0.25846401992455376   0.7820589490422108   0.5828516582565737   0.8349030914844726   0.7163459563685869   0.26818707104558265   0.353680241106759   0.5674790027969111   0.3151479559988224   0.3889985432432684   0.9724260311547991   0.37194363558468974   0.7833905405611205   0.4389387651379187   0.07964567623929604   0.6161937079250903   0.7770714415630412   0.7127197019325895   0.5927511346608791   0.2562035774725487   0.3401613708673031   0.9961468081514423   0.030060142268043558   0.9606281896232727   0.08169735094274931   0.21408785910923145   0.4472084840114699   0.12572509813880012   0.36535139457416244
0.9459007880636489   0.09352824290471089   0.558246095341889   0.05020343857534004   0.5569022448203804   0.1211022117499118   0.18630245975719925   0.26681289801421954   0.11796347968246175   0.041456535510615754   0.570108751832109   0.48974145645117834   0.40524377774987225   0.4487054008497366   0.3139051743595603   0.14958008558387523   0.4090969695984299   0.41864525858169305   0.3532769847362876   0.06788273464112592   0.19500911048919845   0.9714367745702231   0.22755188659748746   0.7025313400669635   0.24910832242554964   0.8779085316655123   0.6693057912555985   0.6523279014916235   0.6922060776051693   0.7568063199156004   0.48300333149839925   0.38551500347740386   0.5742425979227075   0.7153497844049846   0.9128945796662903   0.8957735470262256   0.16899882017283524   0.2666443835552481   0.5989894053067301   0.7461934614423503   0.7599018505744054   0.847999124973555   0.24571242057044243   0.6783107268012244   0.564892740085207   0.8765623504033319   0.018160533972954977   0.9757793867342609   0.3157844176596573   0.9986538187378197   0.3488547427173565   0.32345148524263756   0.6235783400544881   0.2418474988222192   0.8658514112189573   0.9379364817652337   0.04933574213178058   0.5264977144172345   0.952956831552667   0.04216293473900811   0.8803369219589453   0.2598533308619864   0.3539674262459369   0.2959694732966578
0.12043507138453997   0.41185420588843136   0.1082550056754945   0.6176587464954334   0.5555423312993331   0.5352918554850995   0.09009447170253952   0.6418793597611724   0.23975791363967577   0.5366380367472798   0.741239728985183   0.3184278745185349   0.6161795735851877   0.2947905379250606   0.8753883177662258   0.38049139275330124   0.5668438314534071   0.7682928235078261   0.9224314862135589   0.3383284580142931   0.6865069094944618   0.5084394926458397   0.568464059967622   0.04235898471763532   0.5660718381099218   0.09658528675740835   0.4602090542921274   0.42470023822220193   0.010529506810588762   0.5612934312723089   0.3701145825895879   0.7828208784610295   0.770771593170913   0.02465539452502911   0.6288748536044049   0.46439300394249466   0.1545920195857253   0.7298648565999685   0.753486535838179   0.08390161118919344   0.5877481881323182   0.9615720330921425   0.8310550496246203   0.7455731531749004   0.9012412786378564   0.4531325404463027   0.26259098965699834   0.703214168457265   0.33516944052793457   0.35654725368889434   0.8023819353648709   0.27851393023506305   0.32463993371734584   0.7952538224165855   0.43226735277528305   0.4956930517740335   0.5538683405464329   0.7705984278915563   0.8033924991708782   0.03130004783153887   0.39927632096070753   0.040733571291587826   0.04990596333269912   0.9473984366423455
0.8115281328283893   0.07916153819944542   0.21885091370807888   0.20182528346744508   0.9102868541905329   0.6260289977531427   0.9562599240510805   0.4986111150101801   0.5751174136625984   0.26948174406424835   0.1538779886862096   0.220097184775117   0.2504774799452525   0.4742279216476629   0.7216106359109266   0.7244041330010835   0.6966091393988197   0.7036294937561066   0.9182181367400484   0.6931040851695446   0.29733281843811216   0.6628959224645188   0.8683121734073492   0.7457056485271992   0.48580468560972284   0.5837343842650733   0.6494612596992704   0.5438803650597541   0.5755178314191899   0.9577053865119306   0.6932013356481899   0.045269250049574036   0.00040041775659155755   0.6882236424476823   0.5393233469619801   0.825172065274457   0.749922937811339   0.21399572080001933   0.8177127110510536   0.10076793227337354   0.053313798412519355   0.5103662270439128   0.8994945743110052   0.4076638471038289   0.7559809799744072   0.847470304579394   0.03118240090365601   0.6619581985766297   0.2701762943646844   0.2637359203143207   0.38172114120438566   0.11807783351687562   0.6946584629454945   0.3060305338023901   0.6885198055561959   0.07280858346730158   0.6942580451889029   0.6178068913547078   0.14919645859421565   0.24763651819284457   0.9443351073775639   0.40381117055468846   0.331483747543162   0.14686858591947102
0.8910213089650445   0.8934449435107757   0.43198917323215674   0.7392047388156421   0.1350403289906373   0.04597463893138169   0.40080677232850076   0.07724654023901238   0.864864034625953   0.782238718617061   0.019085631124115092   0.9591687067221367   0.1702055716804585   0.4762081848146709   0.33056582556791925   0.8863601232548352   0.4759475264915556   0.8584012934599631   0.18136936697370362   0.6387236050619906   0.5316124191139917   0.4545901229052746   0.8498856194305416   0.49185501914251956   0.6405911101489472   0.5611451793944989   0.41789644619838484   0.7526502803268774   0.50555078115831   0.5151705404631173   0.017089673869884105   0.6754037400878651   0.640686746532357   0.7329318218460562   0.998004042745769   0.7162350333657284   0.4704811748518985   0.2567236370313853   0.6674382171778498   0.8298749101108932   0.9945336483603429   0.3983223435714222   0.48606885020414614   0.19115130504890257   0.4629212292463511   0.9437322206661476   0.6361832307736045   0.699296285906383   0.8223301190974038   0.3825870412716486   0.21828678457521972   0.9466460055795055   0.3167793379390939   0.8674165008085314   0.2011971107053356   0.27124226549164043   0.6760925914067369   0.13448467896247518   0.20319306795956657   0.5550072321259121   0.2056114165548385   0.8777610419310898   0.5357548507817168   0.725132322015019
0.2110777681944956   0.4794386983596677   0.049686000577570666   0.5339810169661163   0.7481565389481445   0.5357064776935201   0.4135027698039661   0.8346847310597334   0.9258264198507407   0.15311943642187148   0.1952159852287464   0.8880387254802279   0.6090470819116467   0.2857029356133401   0.9940188745234108   0.6167964599885875   0.9329544905049098   0.1512182566508649   0.7908258065638443   0.06178922786267533   0.7273430739500713   0.273457214719775   0.2550709557821274   0.3366569058476564   0.5162653057555756   0.7940185163601073   0.20538495520455674   0.80267588888154   0.7681087668074311   0.25831203866658725   0.7918821854005906   0.9679911578218067   0.8422823469566905   0.10519260224471577   0.5966662001718442   0.07995243234157874   0.2332352650450438   0.8194896666313757   0.6026473256484334   0.46315597235299133   0.3002807745401341   0.6682714099805108   0.8118215190845892   0.40136674449031595   0.5729377005900628   0.39481419526073575   0.5567505633024618   0.06470983864265958   0.05667239483448717   0.6007956789006283   0.35136560809790507   0.2620339497611196   0.28856362802705604   0.3424836402340411   0.5594834226973144   0.294042791939313   0.4462812810703655   0.23729103798932533   0.9628172225254702   0.2140903595977342   0.21304601602532172   0.41780137135794965   0.36016989687703677   0.7509343872447429
0.9127652414851877   0.7495299613774389   0.5483483777924476   0.3495676427544269   0.3398275408951249   0.35471576611670314   0.9915978144899859   0.2848578041117673   0.2831551460606377   0.7539200872160747   0.6402322063920808   0.02282385435064776   0.9945915180335817   0.4114364469820337   0.08074878369476633   0.7287810624113348   0.5483102369632161   0.17414540899270833   0.11793156116929614   0.5146907028136006   0.33526422093789443   0.7563440376347587   0.7577616642922593   0.7637563155688577   0.42249897945270676   0.006814076257319829   0.20941328649981178   0.4141886728144308   0.08267143855758186   0.6520983101406167   0.21781547200982598   0.12933086870266342   0.7995162924969441   0.898178222924542   0.5775832656177452   0.10650701435201566   0.8049247744633624   0.4867417759425083   0.4968344819229789   0.37772595194068087   0.25661453750014634   0.3125963669497999   0.37890292075368276   0.8630352491270803   0.9213503165622519   0.5562523293150412   0.6211412564614234   0.09927893355822259   0.49885133710954516   0.5494382530577214   0.41172796996161165   0.6850902607437919   0.4161798985519633   0.8973399429171047   0.19391249795178567   0.5557593920411285   0.6166636060550191   0.9991617199925628   0.6163292323340405   0.44925237768911275   0.8117388315916567   0.5124199440500545   0.11949475041106153   0.07152642574843192
0.5551242940915104   0.19982357710025458   0.7405918296573788   0.20849117662135164   0.6337739775292585   0.6435712477852134   0.11945057319595537   0.10921224306312903   0.1349226404197133   0.09413299472749195   0.7077226032343438   0.4241219823193372   0.71874274186775   0.19679305181038725   0.5138101052825581   0.8683625902782087   0.10207913581273081   0.19763133181782447   0.8974808729485176   0.419110212589096   0.2903403042210741   0.6852113877677699   0.7779861225374561   0.34758378684066404   0.7352160101295637   0.48538781066751535   0.03739429288007735   0.13909261021931243   0.10144203260030525   0.841816562882302   0.917943719684122   0.029880367156183404   0.9665193921805919   0.7476835681548101   0.21022111644977823   0.6057583848368462   0.24777665031284196   0.5508905163444228   0.6964110111672202   0.7373957945586375   0.14569751450011115   0.3532591845265983   0.7989301382187025   0.3182855819695415   0.8553572102790371   0.6680477967588284   0.02094401568124637   0.9707017951288774   0.12014120014947333   0.182659986091313   0.983549722801169   0.8316091849095649   0.01869916754916808   0.340843423209011   0.06560600311704705   0.8017288177533816   0.05217977536857613   0.593159855054201   0.8553848866672688   0.19597043291653535   0.8044031250557342   0.04226933870977822   0.15897387550004866   0.4585746383578979
0.658705610555623   0.6890101541831799   0.36004373728134614   0.1402890563883564   0.8033484002765859   0.02096235742435154   0.33909972160009977   0.169587261259479   0.6832072001271127   0.8383023713330385   0.35554999879893073   0.33797807634991406   0.6645080325779446   0.4974589481240275   0.2899439956818837   0.5362492585965325   0.6123282572093685   0.9042990930698265   0.4345591090146149   0.3402788256799971   0.8079251321536343   0.8620297543600483   0.27558523351456626   0.8817041873220992   0.14921952159801125   0.17301960017686838   0.9155414962332201   0.7414151309337428   0.3458711213214253   0.15205724275251684   0.5764417746331203   0.5718278696742638   0.6626639211943127   0.31375487141947833   0.22089177583418956   0.2338497933243498   0.9981558886163682   0.8162959232954509   0.9309477801523058   0.6976005347278174   0.3858276314069997   0.9119968302256243   0.4963886711376909   0.3573217090478202   0.5779024992533655   0.04996707586557603   0.22080343762312468   0.4756175217257209   0.42868297765535424   0.8769474756887077   0.3052619413899046   0.7342023907919781   0.08281185633392894   0.7248902329361908   0.7288201667567843   0.16237452111771425   0.4201479351396163   0.4111353615167125   0.5079283909225947   0.9285247277933645   0.4219920465232481   0.5948394382212616   0.5769806107702888   0.23092419306554718
0.03616441511624842   0.6828426079956373   0.08059193963259793   0.873602484017727   0.45826191586288295   0.6328755321300613   0.8597885020094732   0.3979849622920061   0.02957893820752871   0.7559280564413536   0.5545265606195687   0.663782571500028   0.9467670818735998   0.03103782350516287   0.8257063938627844   0.5014080503823137   0.5266191467339835   0.6199024619884503   0.3177780029401897   0.5728833225889493   0.10462710021073535   0.02506302376718871   0.7407973921699008   0.3419591295234021   0.06846268509448693   0.3422204157715514   0.6602054525373029   0.4683566455056751   0.6102007692316039   0.7093448836414901   0.8004169505278297   0.07037168321366902   0.5806218310240753   0.9534168272001363   0.24589038990826098   0.40658911171364104   0.6338547491504756   0.9223790036949735   0.42018399604547657   0.9051810613313273   0.10723560241649202   0.3024765417065231   0.10240599310528682   0.33229773874237806   0.0026085022057566773   0.2774135179393344   0.36160860093538594   0.990338609218976   0.9341458171112698   0.9351931021677831   0.701403148398083   0.5219819637133009   0.32394504787966577   0.22584821852629303   0.9009861978702534   0.45161028049963187   0.7433232168555904   0.2724313913261567   0.6550958079619924   0.04502116878599082   0.10946846770511495   0.3500523876311832   0.23491181191651583   0.13984010745466352
0.0022328652886229317   0.04757584592466009   0.13250581881122903   0.8075423687122855   0.9996243630828663   0.7701623279853257   0.7708972178758431   0.8172037594933096   0.06547854597159651   0.8349692258175426   0.06949406947776002   0.2952217957800087   0.7415334980919307   0.6091210072912496   0.16850787160750666   0.8436115152803768   0.9982102812363403   0.336689615965093   0.5134120636455143   0.798590346494386   0.8887418135312253   0.9866372283339098   0.2785002517289984   0.6587502390397225   0.8865089482426024   0.9390613824092497   0.1459944329177694   0.851207870327437   0.8868845851597361   0.168899054423924   0.37509721504192634   0.03400411083412745   0.8214060391881396   0.3339298286063813   0.3056031455641663   0.7387823150541187   0.07987254109620887   0.7248088213151317   0.13709527395665966   0.8951707997737419   0.0816622598598686   0.3881192053500387   0.6236832103111454   0.0965804532793559   0.19292044632864327   0.4014819770161289   0.345182958582147   0.4378302142396334   0.3064114980860409   0.46242059460687923   0.1991885256643776   0.5866223439121964   0.4195269129263048   0.29352154018295523   0.8240913106224513   0.5526182330780689   0.5981208737381651   0.9595917115765739   0.518488165058285   0.8138359180239502   0.5182483326419562   0.23478289026144222   0.38139289110162533   0.9186651182502082
0.43658607278208766   0.8466636849114035   0.75770968079048   0.8220846649708523   0.2436656264534444   0.44518170789527456   0.4125267222083329   0.38425445073121894   0.9372541283674035   0.9827611132883953   0.21333819654395533   0.7976321068190225   0.5177272154410987   0.6892395731054402   0.3892468859215041   0.2450138737409536   0.9196063417029335   0.7296478615288663   0.870758720863219   0.4311779557170034   0.4013580090609773   0.494864971267424   0.48936582976159376   0.5125128374667951   0.9647719362788896   0.6482012863560205   0.7316561489711139   0.6904281724959428   0.7211063098254452   0.20301957846074595   0.3191294267627809   0.30617372176472385   0.7838521814580417   0.22025846517235056   0.10579123021882555   0.5085416149457013   0.266124966016943   0.5310188920669104   0.7165443442973215   0.2635277412047477   0.3465186243140094   0.8013710305380443   0.8457856234341025   0.8323497854877443   0.9451606152530321   0.3065060592706202   0.35641979367250864   0.31983694802094914   0.9803886789741425   0.6583047729145997   0.6247636447013949   0.6294087755250064   0.2592823691486973   0.45528519445385374   0.30563421793861395   0.3232350537602825   0.4754301876906556   0.23502672928150314   0.1998429877197884   0.8146934388145812   0.20930522167371257   0.7040078372145927   0.48329864342246687   0.5511656976098335
0.8627865973597032   0.9026368066765484   0.6375130199883645   0.7188159121220892   0.917625982106671   0.5961307474059283   0.2810932263158558   0.3989789641011401   0.9372373031325285   0.9378259744913287   0.656329581614461   0.7695701885761337   0.6779549339838312   0.4825407800374749   0.350695363675847   0.44633513481585124   0.20252474629317566   0.2475140507559718   0.1508523759560586   0.63164169600127   0.9932195246194631   0.5435062135413791   0.6675537325335917   0.0804759983914365   0.13043292725975994   0.6408694068648306   0.03004071254522725   0.36166008626934726   0.21280694515308893   0.04473865945890233   0.7489474862293715   0.9626811221682072   0.2755696420205604   0.10691268496757368   0.09261790461491048   0.19311093359207346   0.5976147080367292   0.6243719049300988   0.7419225409390635   0.7467757987762222   0.39508996174355354   0.3768578541741269   0.5910701649830048   0.11513410277495223   0.40187043712409043   0.8333516406327478   0.9235164324494132   0.03465810438351573   0.2714375098643305   0.19248223376791718   0.8934757199041858   0.6729980181141685   0.05863056471124158   0.14774357430901483   0.14452823367481443   0.7103168959459613   0.7830609226906812   0.04083088934144116   0.05191032905990395   0.5172059623538878   0.185446214653952   0.41645898441134244   0.3099877881208405   0.7704301635776656
0.7903562529103985   0.039601130237215496   0.7189176231378356   0.6552960608027133   0.38848581578630803   0.20624948960446768   0.7954011906884225   0.6206379564191976   0.11704830592197756   0.01376725583655051   0.9019254707842366   0.9476399383050291   0.058417741210735966   0.8660236815275356   0.7573972371094222   0.23732304235906787   0.2753568185200548   0.8251927921860945   0.7054869080495182   0.72011708000518   0.08991060386610279   0.4087338077747521   0.39549911992867776   0.9496869164275146   0.2995543509557043   0.3691326775375366   0.6765814967908421   0.2943908556248013   0.9110685351693962   0.16288318793306888   0.8811803061024196   0.6737528992056037   0.7940202292474187   0.14911593209651838   0.979254835318183   0.7261129609005745   0.7356024880366827   0.28309225056898274   0.22185759820876083   0.48878991854150666   0.46024566951662793   0.4578994583828882   0.5163706901592426   0.7686728385363266   0.37033506565052515   0.04916565060813614   0.12087157023056484   0.818985922108812   0.07078071469482086   0.6800329730705995   0.4442900734397227   0.5245950664840108   0.1597121795254246   0.5171497851375306   0.5631097673373031   0.8508421672784071   0.3656919502780059   0.36803385304101227   0.5838549320191201   0.12472920637783254   0.6300894622413231   0.08494160247202956   0.3619973338103592   0.6359392878363259
0.1698437927246952   0.6270421440891414   0.8456266436511166   0.8672664492999993   0.79950872707417   0.5778764934810052   0.7247550734205518   0.04828052719118726   0.7287280123793491   0.8978435204104056   0.280464999980829   0.5236854607071765   0.5690158328539245   0.380693735272875   0.717355232643526   0.6728432934287694   0.20332388257591869   0.012659882231862712   0.13350030062440593   0.5481140870509369   0.5732344203345955   0.9277182797598331   0.7715029668140467   0.912174799214611   0.40339062760990035   0.3006761356706918   0.9258763231629301   0.044908349914611706   0.6038819005357303   0.7227996421896866   0.20112124974237838   0.9966278227234244   0.8751538881563812   0.8249561217792809   0.9206562497615494   0.47294236201624795   0.30613805530245664   0.4442623865064059   0.20330101711802337   0.8000990685874786   0.10281417272653795   0.4316025042745432   0.06980071649361744   0.25198498153654175   0.5295797523919424   0.50388422451471   0.2982977496795707   0.3398101823219307   0.12618912478204206   0.20320808884401828   0.37242142651664056   0.29490183240731904   0.5223072242463117   0.4804084466543317   0.17130017677426218   0.2982740096838946   0.6471533360899305   0.6554523248750508   0.2506439270127128   0.8253316476676467   0.3410152807874739   0.21118993836864483   0.04734290989468946   0.025232579080168054
0.23820110806093597   0.7795874340941016   0.9775421934010721   0.7732475975436264   0.7086213556689935   0.27570320957939154   0.6792444437215013   0.4334374152216956   0.5824322308869515   0.07249512073537326   0.30682301720486077   0.13853558281437653   0.06012500664063978   0.5920866740810415   0.13552284043059862   0.8402615731304819   0.41297167055070927   0.9366343492059908   0.8848789134178858   0.014929925462835305   0.07195638976323533   0.725444410837346   0.8375360035231963   0.9896973463826673   0.8337552817022994   0.9458569767432443   0.8599938101221243   0.21644974883904092   0.1251339260333058   0.6701537671638528   0.18074936640062297   0.7830123336173453   0.5427016951463544   0.5976586464284795   0.8739263491957622   0.6444767508029688   0.48257668850571456   0.005571972347438002   0.7384035087651636   0.8042151776724868   0.0696050179550053   0.0689376231414472   0.8535245953472778   0.7892852522096516   0.99764862819177   0.34349321230410124   0.015988591824081487   0.7995879058269844   0.1638933464894706   0.39763623556085687   0.15599478170195719   0.5831381569879434   0.03875942045616479   0.727482468397004   0.9752454153013342   0.800125823370598   0.49605772530981046   0.12982382196852452   0.10131906610557201   0.15564907256762922   0.013481036804095924   0.1242518496210865   0.3629155573404084   0.3514338948951423
0.9438760188490907   0.0553142264796393   0.5093909619931306   0.5621486426854908   0.9462273906573206   0.711821014175538   0.4934023701690491   0.7625607368585064   0.78233404416785   0.31418477861468114   0.3374075884670919   0.17942257987056304   0.7435746237116853   0.586702310217677   0.3621621731657577   0.37929675649996497   0.24751689840187477   0.45687848824915256   0.2608431070601857   0.22364768393233578   0.23403586159777887   0.3326266386280661   0.8979275497197773   0.8722137890371934   0.2901598427486882   0.2773124121484268   0.3885365877266467   0.3100651463517027   0.3439324520913676   0.5654913979728887   0.8951342175575976   0.5475044094931962   0.5615984079235176   0.2513066193582076   0.5577266290905056   0.3680818296226332   0.8180237842118323   0.6646043091405305   0.19556445592474794   0.9887850731226682   0.5705068858099576   0.2077258208913779   0.9347213488645623   0.7651373891903324   0.33647102421217867   0.8750991822633118   0.03679379914478494   0.892923600153139   0.04631118146349042   0.597786770114885   0.6482572114181383   0.5828584538014363   0.7023787293721229   0.03229537214199629   0.7531229938605407   0.035354044308240115   0.14078032144860528   0.7809887527837888   0.19539636477003502   0.6672722146856069   0.322756537236773   0.11638444364325826   0.999831908845287   0.6784871415629388
0.7522496514268154   0.9086586227518804   0.06511055998072487   0.9133497523726064   0.4157786272146368   0.03355944048856858   0.028316760835939935   0.02042615221946738   0.3694674457511464   0.43577267037368356   0.3800595494178017   0.43756769841803106   0.6670887163790236   0.40347729823168726   0.626936555557261   0.40221365410979093   0.5263083949304183   0.6224885454478986   0.43154019078722594   0.734941439424184   0.20355185769364528   0.5061041018046403   0.43170828194193883   0.056454297861245215   0.4513022062668298   0.5974454790527599   0.366597721961214   0.14310454548863885   0.03552357905219301   0.5638860385641913   0.33828096112527406   0.12267839326917146   0.6660561333010466   0.12811336819050775   0.9582214117074723   0.6851106948511404   0.9989674169220231   0.7246360699588205   0.33128485615021136   0.28289704074134947   0.47265902199160476   0.10214752451092195   0.8997446653629854   0.5479556013171655   0.2691071642979595   0.5960434227062816   0.46803638342104653   0.4915013034559203   0.8178049580311296   0.9985979436535217   0.10143866145983256   0.3483967579672814   0.7822813789789367   0.43471190508933044   0.7631577003345585   0.22571836469810996   0.11622524567789001   0.3065985368988227   0.8049362886270861   0.5406076698469695   0.11725782875586696   0.5819624669400022   0.4736514324768748   0.2577106291056201
0.6445988067642622   0.47981494242908024   0.5739067671138894   0.7097550277884546   0.37549164246630273   0.8837715197227985   0.10587038369284285   0.21825372433253432   0.5576866844351731   0.8851735760692768   0.004431722233010293   0.8698569663652529   0.7754053054562364   0.4504616709799463   0.24127402189845176   0.6441386016671429   0.6591800597783464   0.14386313408112364   0.4363377332713656   0.10353093182017337   0.5419222310224795   0.5619006671411214   0.9626863007944908   0.8458203027145533   0.8973234242582172   0.08208572471204122   0.3887795336806014   0.1360652749260987   0.5218317817919146   0.19831420498924265   0.28290914998775857   0.9178115505935645   0.9641450973567415   0.31314062891996586   0.27847742775474826   0.04795458422831153   0.18873979190050505   0.8626789579400195   0.0372034058562965   0.40381598256116863   0.5295597321221587   0.7188158238588959   0.6008656725849308   0.30028505074099526   0.9876375010996792   0.1569151567177744   0.63817937179044   0.45446474802644193   0.09031407684146195   0.07482943200573319   0.24939983810983865   0.3183994731003432   0.5684822950495474   0.8765152270164905   0.96649068812208   0.4005879225067788   0.6043371976928059   0.5633745980965247   0.6880132603673318   0.3526333382784673   0.41559740579230087   0.7006956401565052   0.6508098545110353   0.9488173557172987
0.8860376736701422   0.9818798162976093   0.04994418192610441   0.6485323049763034   0.898400172570463   0.8249646595798349   0.41176481013566435   0.1940675569498615   0.808086095729001   0.7501352275741018   0.1623649720258257   0.8756680838495182   0.23960380067945367   0.8736200005576112   0.19587428390374564   0.4750801613427394   0.6352666029866477   0.3102454024610865   0.5078610235364138   0.1224468230642721   0.21966919719434685   0.6095497623045812   0.8570511690253786   0.1736294673469734   0.3336315235242046   0.627669946006972   0.8071069870992742   0.52509716237067   0.43523135095374155   0.802705286427137   0.3953421769636098   0.33102960542080845   0.6271452552247405   0.05257005885303529   0.2329772049377841   0.45536152157129023   0.3875414545452868   0.1789500582954241   0.03710292103403844   0.9802813602285508   0.752274851558639   0.8687046558343376   0.5292418974976246   0.8578345371642787   0.5326056543642922   0.2591548935297563   0.672190728472246   0.6842050698173053   0.19897413084008764   0.6314849475227844   0.8650837413729718   0.15910790744663536   0.7637427798863461   0.8287796610956473   0.4697415644093621   0.8280783020258269   0.13659752466160557   0.776209602242612   0.236764359471578   0.37271678045453666   0.7490560701163187   0.5972595439471879   0.19966143843753956   0.3924354202259859
0.9967812185576796   0.7285548881128503   0.670419540939915   0.5346008830617072   0.4641755641933874   0.469399994583094   0.9982288124676689   0.8503958132444018   0.2652014333532998   0.8379150470603096   0.13314507109469703   0.6912879057977666   0.5014586534669537   0.00913538596466235   0.663403506685335   0.8632096037719397   0.3648611288053482   0.23292578372205033   0.42663914721375695   0.49049282331740296   0.6158050586890295   0.6356662397748624   0.22697770877621737   0.09805740309141708   0.6190238401313498   0.9071113516620121   0.5565581678363024   0.5634565200297099   0.15484827593796235   0.43771135707891806   0.5583293553686335   0.713060706785308   0.8896468425846625   0.5997963100186084   0.4251842842739364   0.021772800987541484   0.3881881891177088   0.5906609240539461   0.7617807775886015   0.15856319721560183   0.023327060312360613   0.35773514033189574   0.3351416303748445   0.6680703738981989   0.4075220016233312   0.7220689005570333   0.10816392159862714   0.5700129708067818   0.7884981614919814   0.8149575488950213   0.5516057537623248   0.006556450777071891   0.633649885554019   0.3772461918161032   0.9932763983936913   0.29349574399176387   0.7440030429693565   0.7774498817974947   0.5680921141197549   0.2717229430042224   0.3558148538516477   0.1867889577435487   0.8063113365311534   0.11315974578862055
0.3324877935392871   0.829053817411653   0.4711697061563089   0.4450893718904217   0.9249657919159558   0.10698491685461964   0.36300578455768173   0.8750764010836399   0.1364676304239745   0.2920273679595984   0.8114000307953569   0.868519950306568   0.5028177448699555   0.9147811761434952   0.8181236324016657   0.5750242063148041   0.758814701900599   0.13733129434600044   0.25003151828191084   0.3033012633105817   0.4029998480489513   0.9505423366024518   0.44372018175075745   0.19014151752196118   0.07051205450966425   0.12148851919079878   0.9725504755944485   0.7450521456315395   0.14554626259370834   0.014503602336179146   0.6095446910367668   0.8699757445478996   0.009078632169733846   0.7224762343765808   0.7981446602414098   0.0014557942413316396   0.5062608872997784   0.8076950582330855   0.9800210278397441   0.4264315879265275   0.7474461853991794   0.6703637638870851   0.7299895095578334   0.1231303246159458   0.34444633735022806   0.7198214272846334   0.2862693278070759   0.9329888070939846   0.2739342828405638   0.5983329080938345   0.31371885221262735   0.18793666146244511   0.1283880202468555   0.5838293057576555   0.7041741611758605   0.3179609169145455   0.11930938807712164   0.8613530713810746   0.9060295009344507   0.31650512267321385   0.6130485007773433   0.053658013147989125   0.9260084730947066   0.8900735347466863
0.8656023153781639   0.383294249260904   0.19601896353687323   0.7669432101307405   0.5211559780279358   0.6634728219762707   0.9097496357297974   0.8339544030367559   0.24722169518737194   0.06513991388243606   0.59603078351717   0.6460177415743108   0.11883367494051647   0.4813106081247806   0.8918566223413095   0.3280568246597653   0.9995242868633948   0.6199575367437059   0.9858271214068587   0.01155170198655149   0.38647578608605154   0.5662995235957168   0.05981864831215217   0.12147816723986518   0.5208734707078877   0.1830052743348128   0.8637996847752789   0.35453495710912464   0.9997174926799519   0.5195324523585422   0.9540500490454816   0.5205805540723688   0.7524957974925799   0.4543925384761061   0.3580192655283116   0.874562812498058   0.6336621225520634   0.9730819303513255   0.4661626431870022   0.5465059878382926   0.6341378356886687   0.35312439360761955   0.48033552178014344   0.5349542858517411   0.2476620496026171   0.7868248700119027   0.42051687346799127   0.41347611861187594   0.7267885788947294   0.60381959567709   0.5567171886927124   0.05894116150275129   0.7270710862147775   0.08428714331854778   0.6026671396472307   0.5383606074303825   0.9745752887221976   0.6298946048424416   0.24464787411891917   0.6637977949323246   0.34091316617013406   0.6568126744911162   0.778485230931917   0.11729180709403196
0.7067753304814655   0.30368828088349664   0.2981497091517735   0.5823375212422909   0.45911328087884834   0.5168634108715939   0.8776328356837823   0.16886140263041488   0.7323247019841189   0.913043815194504   0.3209156469910699   0.10992024112766358   0.005253615769341463   0.8287566718759563   0.718248507343839   0.571559633697281   0.0306783270471439   0.19886206703351453   0.47360063322491996   0.9077618387649564   0.6897651608770098   0.5420493925423983   0.695115402293003   0.7904700316709244   0.9829898303955443   0.23836111165890164   0.3969656931412295   0.20813251042863365   0.523876549516696   0.7214977007873077   0.5193328574574472   0.03927110779821879   0.791551847532577   0.8084538855928037   0.19841721046637736   0.9293508666705552   0.7862982317632355   0.9796972137168475   0.48016870312253823   0.3577912329732742   0.7556199047160916   0.780835146683333   0.006568069897618301   0.4500293942083177   0.06585474383908188   0.2387857541409347   0.3114526676046153   0.6595593625373932   0.0828649134435375   0.00042464248203305825   0.9144869744633859   0.45142685210875955   0.5589883639268415   0.2789269416947253   0.39515411700593867   0.4121557443105408   0.7674365163942645   0.4704730561019216   0.1967369065395613   0.4828048776399856   0.9811382846310288   0.4907758423850741   0.716568203417023   0.1250136446667114
0.22551837991493714   0.7099406957017411   0.7100001335194047   0.6749842504583937   0.15966363607585526   0.47115494156080634   0.3985474659147894   0.015424887921000439   0.07679872263231777   0.4707302990787733   0.48406049145140356   0.5639980358122408   0.5178103587054763   0.19180335738404797   0.0889063744454649   0.1518422915017001   0.7503738423112118   0.7213303012821264   0.8921694679059036   0.6690374138617146   0.769235557680183   0.23055445889705228   0.17560126448888055   0.5440237691950032   0.5437171777652459   0.5206137631953112   0.4656011309694758   0.8690395187366095   0.3840535416893906   0.049458821634504845   0.0670536650546864   0.853614630815609   0.30725481905707286   0.5787285225557316   0.5829931736032828   0.2896165950033681   0.7894444603515965   0.38692516517168357   0.49408679915781795   0.13777430350166806   0.039070618040384676   0.6655948638895572   0.6019173312519144   0.4687368896399535   0.26983506036020166   0.43504040499250496   0.4263160667630338   0.9247131204449505   0.7261178825949558   0.9144266417971937   0.9607149357935579   0.05567360170834097   0.34206434090556515   0.8649678201626889   0.8936612707388716   0.20205897089273198   0.034809521848492335   0.2862392976069573   0.3106680971355887   0.9124423758893638   0.2453650614968958   0.8993141324352738   0.8165812979777707   0.7746680723876957
0.20629444345651113   0.23371926854571654   0.21466396672585636   0.3059311827477422   0.9364593830963095   0.7986788635532116   0.7883478999628226   0.3812180623027918   0.2103415005013537   0.8842522217560179   0.8276329641692646   0.32554446059445086   0.8682771595957886   0.019284401593329024   0.933971693430393   0.12348548970171888   0.8334676377472962   0.7330451039863717   0.6233035962948044   0.21104311381235505   0.5881025762504004   0.833730971551098   0.8067222983170337   0.43637504142465927   0.38180813279388925   0.6000117030053814   0.5920583315911773   0.13044385867691705   0.4453487496975798   0.8013328394521698   0.8037104316283548   0.7492257963741252   0.23500724919622612   0.9170806176961519   0.9760774674590901   0.4236813357796744   0.36673008960043757   0.8977962161028229   0.04210577402869708   0.3001958460779555   0.5332624518531414   0.16475111211645116   0.4188021777338927   0.08915273226560046   0.945159875602741   0.3310201405653532   0.612079879416859   0.6527776908409412   0.5633517428088517   0.7310084375599718   0.020021547825681805   0.5223338321640241   0.11800299311127192   0.9296755981078021   0.2163111161973271   0.7731080357898988   0.8829957439150458   0.012594980411650192   0.24023364873823697   0.34942670001022447   0.5162656543146082   0.11479876430882734   0.19812787470953988   0.04923085393226897
0.9830032024614668   0.9500476521923762   0.7793256969756471   0.9600781216666685   0.03784332685872581   0.619027511627023   0.1672458175587881   0.30730043082572733   0.47449158404987407   0.8880190740670512   0.14722426973310626   0.7849665986617033   0.35648859093860213   0.9583434759592491   0.9309131535357792   0.011858562871804326   0.4734928470235564   0.9457484955475989   0.6906795047975423   0.6624318628615798   0.9572271927089482   0.8309497312387715   0.49255163008800235   0.6132010089293108   0.9742239902474813   0.8809020790463953   0.7132259331123552   0.6531228872626423   0.9363806633887555   0.2618745674193724   0.5459801155535671   0.34582245643691506   0.46188907933888146   0.37385549335232127   0.3987558458204608   0.5608558577752119   0.10540048840027928   0.4155120173930722   0.4678426922846816   0.5489972949034075   0.631907641376723   0.4697635218454734   0.7771631874871394   0.8865654320418277   0.6746804486677748   0.6388137906067018   0.28461155739913707   0.2733644231125168   0.7004564584202935   0.7579117115603066   0.5713856242867819   0.6202415358498744   0.764075795031538   0.49603714414093414   0.02540550873321482   0.2744190794129594   0.3021867156926565   0.12218165078861287   0.626649662912754   0.7135632216377475   0.1967862272923772   0.7066696333955407   0.15880697062807236   0.16456592673434003
0.5648785859156543   0.23690611155006727   0.38164378314093295   0.27800049469251237   0.8901981372478794   0.5980923209433654   0.09703222574179587   0.004636071579995597   0.18974167882758602   0.8401806093830589   0.525646601455014   0.38439453573012117   0.4256658837960481   0.34414346524212475   0.5002410927217992   0.1099754563171618   0.12347916810339157   0.2219618144535119   0.8735914298090451   0.3964122346794143   0.9266929408110144   0.5152921810579713   0.7147844591809728   0.23184630794507421   0.36181435489536007   0.27838606950790395   0.33314067604003983   0.9538458132525618   0.4716162176474806   0.6802937485645385   0.23610845029824395   0.9492097416725662   0.28187453881989455   0.8401131391814797   0.7104618488432299   0.564815205942445   0.8562086550238465   0.49596967393935487   0.21022075612143085   0.45483974962528323   0.7327294869204549   0.274007859485843   0.33662932631238573   0.058427514945868994   0.8060365461094405   0.7587156784278717   0.621844867131413   0.8265812070007947   0.44422219121408046   0.48032960891996773   0.28870419109137313   0.872735393748233   0.9726059735666   0.8000358603554292   0.052595740793129175   0.9235256520756667   0.6907314347467054   0.9599227211739496   0.3421338919498992   0.35871044613322167   0.8345227797228589   0.4639530472345947   0.13191313582846834   0.9038706965079384
0.101793292802404   0.18994518774875171   0.7952838095160826   0.8454431815620694   0.2957567466929635   0.43122950932088   0.1734389423846697   0.018861974561274662   0.851534555478883   0.9508999004009122   0.8847347512932966   0.1461265808130417   0.8789285819122831   0.150864040045483   0.8321390105001674   0.22260092873737497   0.1881971471655777   0.19094131887153346   0.4900051185502682   0.8638904826041532   0.3536743674427188   0.7269882716369388   0.3580919827217999   0.9600197860962149   0.2518810746403148   0.537043083888187   0.5628081732057172   0.11457660453414538   0.9561243279473514   0.10581357456730701   0.3893692308210476   0.09571462997287072   0.10458977246846836   0.1549136741663948   0.504634479527751   0.949588049159829   0.2256611905561853   0.004049634120911755   0.6724954690275836   0.7269871204224541   0.037464043390607604   0.8131083152493783   0.18249035047731538   0.8630966378183008   0.6837896759478889   0.08612004361243956   0.8243983677555156   0.903076851722086   0.431908601307574   0.5490769597242525   0.26159019454979826   0.7885002471879405   0.47578427336022266   0.4432633851569455   0.8722209637287507   0.6927856172150698   0.3711945008917543   0.28834971099055073   0.36758648420099976   0.7431975680552408   0.14553331033556902   0.284300076869639   0.6950910151734162   0.01621044763278677
0.10806926694496141   0.47119176162026066   0.5126006646961008   0.15311380981448597   0.42427959099707263   0.38507171800782114   0.6882022969405853   0.2500369580924   0.9923709896894986   0.8359947582835686   0.426612102390787   0.46153671090445947   0.5165867163292759   0.39273137312662304   0.5543911386620363   0.7687510936893895   0.1453922154375216   0.10438166213607229   0.1868046544610365   0.025553525634148755   0.9998589051019525   0.8200815852664333   0.49171363928762035   0.009343078001361985   0.8917896381569912   0.3488898236461726   0.9791129745915196   0.856229268186876   0.46751004715991856   0.9638181056383515   0.29091067765093426   0.6061923100944759   0.47513905747041996   0.1278233473547829   0.8642985752601473   0.14465559919001653   0.9585523411411441   0.7350919742281599   0.30990743659811104   0.37590450550062693   0.8131601257036225   0.6307103120920876   0.12310278213707451   0.3503509798664782   0.8133012206016699   0.8106287268256542   0.6313891428494541   0.3410079018651162   0.9215115824446788   0.4617389031794817   0.6522761682579347   0.4847786336782402   0.45400153528476017   0.49792079754113017   0.36136549060700035   0.8785863235837642   0.9788624778143402   0.37009745018634727   0.49706691534685304   0.7339307243937477   0.02031013667319618   0.6350054759581873   0.187159478748742   0.35802621889312075
0.20715001096957372   0.0042951638660998145   0.0640566966116675   0.007675239026642556   0.3938487903679038   0.19366643704044553   0.43266755376221333   0.6666673371615264   0.4723372079232251   0.7319275338609639   0.7803913855042788   0.18188870348328615   0.01833567263846487   0.2340067363198337   0.41902589489727843   0.3033023798995219   0.03947319482412463   0.8639092861334865   0.9219589795504254   0.5693716555057742   0.019163058150928454   0.22890381017529907   0.7347995008016833   0.21134543661265348   0.8120130471813547   0.22460864630919924   0.6707428041900159   0.20367019758601093   0.41816425681345093   0.030942209268753705   0.2380752504278025   0.5370028604244845   0.9458270488902258   0.2990146754077898   0.45768386492352375   0.3551141569411984   0.927491376251761   0.06500793908795612   0.03865797002624537   0.05181177704167651   0.8880181814276363   0.20109865295446966   0.11669899047582   0.48244012153590227   0.8688551232767079   0.9721948427791706   0.38189948967413667   0.2710946849232488   0.05684207609535317   0.7475861964699714   0.7111566854841208   0.06742448733723787   0.6386778192819023   0.7166439872012177   0.4730814350563183   0.5304216269127533   0.6928507703916764   0.4176293117934278   0.015397570132794514   0.17530746997155486   0.7653593941399154   0.3526213727054717   0.9767396001065491   0.12349569292987835
0.877341212712279   0.15152271975100204   0.8600406096307291   0.6410555713939761   0.008486089435571104   0.17932787697183145   0.4781411199565925   0.3699608864707273   0.951644013340218   0.43174168050186007   0.7669844344724717   0.3025363991334894   0.3129661940583157   0.7150976933006424   0.2939029994161534   0.7721147722207361   0.6201154236666393   0.2974683815072146   0.27850542928335886   0.5968073022491812   0.8547560295267239   0.9448470088017429   0.3017658291768097   0.4733116093193029   0.9774148168144449   0.7933242890507408   0.4417252195460806   0.8322560379253268   0.9689287273788738   0.6139964120789094   0.9635840995894881   0.46229515145459954   0.017284714038655884   0.18225473157704933   0.1965996651170164   0.15975875232111017   0.7043185199803402   0.4671570382764069   0.902696665700863   0.3876439801003741   0.08420309631370088   0.16968865676919234   0.6241912364175041   0.7908366778511928   0.22944706678697693   0.22484164796744946   0.32242540724069435   0.31752506853188994   0.25203224997253204   0.4315173589167086   0.8807001876946138   0.4852690306065631   0.28310352259365823   0.8175209468377992   0.9171160881051257   0.022973879151963597   0.26581880855500234   0.6352662152607499   0.7205164229881093   0.8632151268308534   0.5615002885746622   0.16810917698434297   0.8178197572872462   0.47557114673047934
0.47729719226096123   0.9984205202151506   0.19362852086974214   0.6847344688792865   0.24785012547398433   0.7735788722477012   0.8712031136290478   0.3672094003473966   0.9958178755014523   0.34206151333099255   0.990502925934434   0.8819403697408335   0.7127143529077941   0.5245405664931934   0.07338683782930831   0.8589664905888698   0.4468955443527918   0.8892743512324435   0.3528704148411991   0.9957513637580163   0.8853952557781296   0.7211651742481006   0.5350506575539528   0.520180217027537   0.4080980635171684   0.7227446540329499   0.3414221366842107   0.8354457481482505   0.16024793804318405   0.9491657817852487   0.4702190230551629   0.46823634780085394   0.16443006254173176   0.6071042684542561   0.47971609712072893   0.5862959780600205   0.45171570963393765   0.08256370196106279   0.4063292592914206   0.7273294874711508   0.004820165281145913   0.19328935072861933   0.05345884445022156   0.7315781237131344   0.11942490950301629   0.4721241764805188   0.5184081868962688   0.21139790668559738   0.7113268459858479   0.7493795224475689   0.1769860502120581   0.37595215853734687   0.5510789079426639   0.8002137406623202   0.7067670271568952   0.9077158107364929   0.38664884540093214   0.19310947220806407   0.22705093003616625   0.3214198326764724   0.9349331357669944   0.11054577024700128   0.8207216707447457   0.5940903452053217
0.9301129704858485   0.917256419518382   0.7672628262945241   0.8625122214921872   0.8106880609828323   0.44513224303786314   0.24885463939825533   0.6511143148065899   0.09936121499698432   0.6957527205902942   0.07186858918619723   0.275162156269243   0.5482823070543205   0.895538979927974   0.36510156202930205   0.3674463455327501   0.1616334616533883   0.70242950771991   0.1380506319931358   0.0460265128562777   0.22670032588639386   0.5918837374729087   0.31732896124839016   0.45193616765095607   0.2965873554005453   0.6746273179545267   0.550066134953866   0.5894239461587688   0.485899294417713   0.22949507491666354   0.3012114955556107   0.9383096313521789   0.3865380794207287   0.5337423543263693   0.2293429063694135   0.6631474750829359   0.8382557723664082   0.6382033743983953   0.8642413443401115   0.2957011295501859   0.6766223107130199   0.9357738666784853   0.7261907123469756   0.24967461669390817   0.44992198482662615   0.34389012920557666   0.4088617510985855   0.7977384490429521   0.15333462942608084   0.6692628112510499   0.8587956161447194   0.2083145028841833   0.6674353350083678   0.4397677363343864   0.5575841205891087   0.2700048715320043   0.28089725558763906   0.9060253820080171   0.3282412142196952   0.6068573964490683   0.4426414832212308   0.2678220076096219   0.46399986987958375   0.3111562668988825
0.7660191725082108   0.33204814093113655   0.7378091575326081   0.06148165020497433   0.31609718768158473   0.98815801172556   0.32894740643402254   0.2637432011620222   0.16276255825550387   0.31889520047451   0.4701517902893031   0.05542869827783893   0.4953272232471361   0.8791274641401235   0.9125676697001943   0.7854238267458346   0.214429967659497   0.9731020821321065   0.5843264554804991   0.17856643029676622   0.7717884844382662   0.7052800745224845   0.1203265856009154   0.8674101633978837   0.005769311930055356   0.373231933591348   0.38251742806830735   0.8059285131929094   0.6896721242484707   0.3850739218657881   0.05357002163428479   0.5421853120308872   0.5269095659929668   0.06617872139127814   0.5834182313449817   0.48675661375304824   0.03158234274583068   0.1870512572511546   0.6708505616447873   0.7013327870072136   0.8171523750863336   0.21394917511904818   0.0865241061642882   0.5227663567104474   0.045363890648067486   0.5086691005965636   0.9661975205633728   0.6553561933125637   0.039594578718012134   0.1354371670052156   0.5836800924950655   0.8494276801196543   0.3499224544695415   0.7503632451394275   0.5301100708607807   0.30724236808876715   0.8230128884765747   0.6841845237481494   0.9466918395157989   0.8204857543357189   0.791430545730744   0.4971332664969948   0.27584127787101165   0.11915296732850533
0.9742781706444104   0.2831840913779466   0.18931717170672344   0.5963866106180579   0.9289142799963429   0.774514990781383   0.22311965114335064   0.9410304173054942   0.8893197012783307   0.6390778237761674   0.6394395586482852   0.09160273718583989   0.5393972468087892   0.8887145786367399   0.1093294877875045   0.7843603690970727   0.7163843583322145   0.2045300548885905   0.16263764827170551   0.9638746147613537   0.9249538126014705   0.7073967883915957   0.8867963704006939   0.8447216474328484   0.9506756419570601   0.4242126970136491   0.6974791986939705   0.2483350368147905   0.021761361960717266   0.6496977062322662   0.4743595475506198   0.3073046195092963   0.13244166068238653   0.01061988245609876   0.8349199889023347   0.2157018823234564   0.5930444138735973   0.12190530381935889   0.7255905011148301   0.4313415132263837   0.8766600555413827   0.9173752489307684   0.5629528528431247   0.4674668984650299   0.9517062429399122   0.20997846053917266   0.6761564824424308   0.6227452510321815   0.0010306009828521462   0.7857657635255235   0.9786772837484603   0.374410214217391   0.9792692390221349   0.13606805729325738   0.5043177361978405   0.06710559470809473   0.8468275783397483   0.12544817483715864   0.6693977472955058   0.8514037123846383   0.25378316446615107   0.0035428710177997464   0.9438072461806757   0.4200621991582546
0.3771231089247683   0.08616762208703135   0.3808543933375511   0.9525953006932246   0.425416865984856   0.8761891615478586   0.7046979108951203   0.32985004966104314   0.4243862650020039   0.09042339802233516   0.72602062714666   0.9554398354436521   0.44511702597986896   0.9543553407290778   0.22170289094881954   0.8883342407355574   0.5982894476401206   0.8289071658919192   0.5523051436533136   0.03693052835091908   0.3445062831739696   0.8253642948741193   0.6084978974726379   0.6168683291926644   0.9673831742492013   0.739196672787088   0.22764350413508685   0.6642730284994398   0.5419663082643453   0.8630075112392294   0.5229455932399665   0.33442297883839667   0.11758004326234141   0.7725841132168941   0.7969249660933064   0.37898314339474454   0.6724630172824724   0.8182287724878164   0.575222075144487   0.49064890265918715   0.07417356964235178   0.9893216065958973   0.022916931491173274   0.45371837430826806   0.7296672864683822   0.16395731172177788   0.4144190340185353   0.8368500451156036   0.7622841122191809   0.42476063893468985   0.18677552988344845   0.17257701661616376   0.22031780395483563   0.5617531276954606   0.6638299366434819   0.8381540377777671   0.10273776069249421   0.7891690144785664   0.8669049705501755   0.4591708943830226   0.4302747434100218   0.97094024199075   0.29168289540568854   0.9685219917238355
0.35610117376767003   0.9816186353948527   0.26876596391451524   0.5148036174155675   0.6264338872992878   0.8176613236730748   0.8543469298959799   0.6779535722999639   0.8641497750801069   0.39290068473838496   0.6675714000125315   0.5053765556838   0.6438319711252714   0.8311475570429244   0.003741463369049507   0.6672225179060329   0.5410942104327771   0.04197854256435801   0.13683649281887406   0.20805162352301038   0.11081946702275527   0.07103830057360803   0.8451535974131855   0.2395296317991749   0.7547182932550852   0.08941966517875534   0.5763876334986703   0.7247260143836075   0.12828440595579743   0.2717583415056805   0.7220407036026903   0.04677244208364366   0.2641346308756905   0.8788576567672955   0.05446930359015894   0.5413958863998436   0.6203026597504192   0.04771009972437119   0.05072784022110943   0.8741733684938107   0.07920844931764212   0.005731557160013173   0.9138913474022354   0.6661217449708002   0.9683889822948868   0.9346932565864051   0.06873774998904984   0.4265921131716253   0.21367068903980158   0.8452735914076498   0.4923501164903795   0.7018660987880179   0.08538628308400416   0.5735152499019692   0.7703094128876892   0.6550936567043741   0.8212516522083136   0.6946575931346737   0.7158401092975302   0.1136977703045306   0.20094899245789444   0.6469474934103026   0.6651122690764207   0.23952440181071996
0.12174054314025233   0.6412159362502894   0.7512209216741854   0.5734026568399198   0.1533515608453655   0.7065226796638842   0.6824831716851355   0.14681054366829438   0.9396808718055639   0.8612490882562344   0.190133055194756   0.44494444488027657   0.8542945887215597   0.28773383835426514   0.41982364230706687   0.7898507881759024   0.0330429365132461   0.5930762452195915   0.7039835330095366   0.6761530178713717   0.8320939440553516   0.9461287518092889   0.038871263933115865   0.4366286160606518   0.7103534009150994   0.3049128155589996   0.2876503422589305   0.8632259592207321   0.5570018400697339   0.5983901358951154   0.6051671705737949   0.7164154155524377   0.6173209682641699   0.737141047638881   0.4150341153790389   0.27147097067216114   0.7630263795426102   0.44940720928461586   0.9952104730719721   0.48162018249625876   0.7299834430293641   0.8563309640650244   0.29122694006243544   0.805467164624887   0.8978894989740124   0.9102022122557355   0.25235567612931953   0.3688385485642352   0.1875360980589131   0.605289396696736   0.964705333870389   0.5056125893435032   0.6305342579891793   0.006899260801620546   0.35953816329659416   0.7891971737910655   0.013213289725009328   0.26975821316273957   0.9445040479175553   0.5177262031189043   0.25018691018239914   0.8203510038781237   0.9492935748455832   0.03610602062264551
0.520203467153035   0.9640200398130992   0.6580666347831478   0.2306388559977585   0.6223139681790226   0.05381782755736368   0.4057109586538282   0.8618003074335233   0.4347778701201095   0.44852843086062777   0.4410056247834392   0.3561877180900202   0.8042436121309302   0.4416291700590072   0.08146746148684501   0.5669905442989548   0.791030322405921   0.17187095689626763   0.13696341356928976   0.049264341180050464   0.5408434122235217   0.351519953018144   0.18766983872370654   0.013158320557404955   0.020639945070486724   0.3874999132050448   0.5296032039405587   0.7825194645596465   0.3983259768914641   0.3336820856476811   0.1238922452867305   0.9207191571261232   0.9635481067713546   0.8851536547870533   0.6828866205032913   0.564531439036103   0.15930449464042434   0.4435244847280462   0.6014191590164463   0.9975408947371482   0.3682741722345034   0.2716535278317785   0.46445574544715656   0.9482765535570977   0.8274307600109816   0.9201335748136346   0.27678590672345005   0.9351182329996929   0.8067908149404949   0.5326336616085897   0.7471827027828912   0.15259876844004636   0.40846483804903083   0.19895157596090868   0.6232904574961607   0.2318796113139232   0.4449167312776762   0.3137979211738553   0.9404038369928694   0.6673481722778202   0.2856122366372519   0.8702734364458091   0.3389846779764231   0.669807277540672
0.9173380644027485   0.5986199086140307   0.8745289325292666   0.7215307239835742   0.08990730439176685   0.6784863338003961   0.5977430258058165   0.7864124909838814   0.28311648945127194   0.1458526721918064   0.8505603230229253   0.6338137225438351   0.8746516514022411   0.9469010962308977   0.22726986552676448   0.4019341112299118   0.4297349201245649   0.6331031750570424   0.28686602853389503   0.7345859389520916   0.14412268348731302   0.7628297386112333   0.9478813505574719   0.0647786614114196   0.22678461908456454   0.16420982999720257   0.07335241802820539   0.3432479374278454   0.13687731469279768   0.4857234961968064   0.47560939222238885   0.556835446443964   0.8537608252415257   0.339870824005   0.6250490691994636   0.9230217239001289   0.9791091738392846   0.3929697277741023   0.39777920367269914   0.5210876126702172   0.5493742537147197   0.7598665527170598   0.11091317513880411   0.7865016737181256   0.4052515702274067   0.9970368141058266   0.16303182458133217   0.721723012306706   0.17846695114284217   0.832826984108624   0.08967940655312678   0.3784750748788606   0.04158963645004449   0.3471034879118176   0.6140700143307379   0.8216396284348966   0.18782881120851874   0.007232663906817637   0.9890209451312743   0.8986179045347676   0.2087196373692341   0.6142629361327153   0.5912417414585751   0.3775302918645505
0.6593453836545143   0.8543963834156555   0.48032856631977106   0.5910286181464249   0.2540938134271077   0.8573595693098289   0.31729674173843886   0.8693056058397189   0.07562686228426549   0.024532585201204878   0.22761733518531208   0.49083053096085827   0.034037225834221   0.6774290972893873   0.6135473208545742   0.6691909025259617   0.8462084146257023   0.6701964333825696   0.6245263757232998   0.770572997991194   0.6374887772564681   0.05593349724985423   0.03328463426472471   0.3930427061266435   0.9781433936019538   0.2015371138341987   0.5529560679449537   0.8020140879802187   0.7240495801748461   0.34417754452436977   0.23565932620651478   0.9327084821404997   0.6484227178905806   0.3196449593231649   0.008041991021202708   0.44187795117964146   0.6143854920563596   0.6422158620337777   0.39449467016662854   0.7726870486536798   0.7681770774306573   0.972019428651208   0.7699682944433287   0.0021140506624857877   0.1306883001741892   0.9160859314013539   0.736683660178604   0.6090713445358422   0.1525449065722354   0.7145488175671552   0.18372759223365032   0.8070572565556237   0.4284953263973893   0.37037127304278533   0.9480682660271356   0.8743487744151239   0.7800726085068087   0.050726313719620435   0.9400262750059328   0.43247082323548247   0.16568711645044906   0.40851045168584277   0.5455316048393043   0.6597837745818027
0.3975100390197917   0.4364910230346347   0.7755633103959756   0.6576697239193169   0.2668217388456025   0.5204050916332809   0.03887965021737161   0.04859837938347463   0.11427683227336709   0.8058562740661258   0.8551520579837213   0.24154112282785098   0.6857815058759777   0.4354850010233405   0.9070837919565857   0.3671923484127271   0.9057088973691692   0.38475868730372004   0.967057516950653   0.9347215251772446   0.7400217809187201   0.9762482356178772   0.4215259121113487   0.2749377505954419   0.34251174189892836   0.5397572125832425   0.6459626017153731   0.617268026676125   0.07569000305332584   0.019352120949961596   0.6070829514980015   0.5686696472926503   0.9614131707799587   0.2134958468838358   0.7519308935142802   0.32712852446479934   0.27563166490398094   0.7780108458604954   0.8448471015576944   0.9599361760520723   0.36992276753481185   0.3932521585567753   0.8777895846070415   0.02521465087482773   0.6299009866160918   0.4170039229388981   0.4562636724956928   0.7502769002793859   0.2873892447171635   0.8772467103556556   0.8103010707803197   0.13300887360326086   0.21169924166383763   0.857894589405694   0.20321811928231814   0.5643392263106105   0.2502860708838789   0.6443987425218582   0.4512872257680379   0.23721070184581114   0.9746544059798979   0.8663878966613628   0.6064401242103435   0.27727452579373885
0.6047316384450862   0.47313573810458753   0.7286505396033021   0.2520598749189111   0.9748306518289943   0.05613181516568941   0.27238686710760923   0.5017829746395253   0.6874414071118309   0.1788851048100338   0.4620857963272896   0.3687741010362644   0.47574216544799325   0.3209905154043398   0.25886767704497143   0.8044348747256539   0.22545609456411433   0.6765917728824816   0.8075804512769335   0.5672241728798427   0.25080168858421636   0.8102038762211188   0.20114032706659   0.28994964708610393   0.6460700501391303   0.33706813811653125   0.47248978746328796   0.03788977216719282   0.671239398310136   0.28093632295084187   0.2001029203556787   0.5361067975276675   0.9837979911983051   0.10205121814080806   0.7380171240283891   0.16733269649140317   0.5080558257503119   0.7810607027364682   0.47914944698341766   0.36289782176574925   0.2825997311861976   0.10446892985398662   0.6715689957064842   0.7956736488859065   0.03179804260198119   0.29426505363286787   0.4704286686398942   0.5057240017998026   0.3857279924628509   0.9571969155163366   0.9979388811766062   0.4678342296326098   0.7144885941527149   0.6762605925654948   0.7978359608209274   0.9317274321049422   0.7306906029544098   0.5742093744246867   0.05981883679253838   0.7643947356135391   0.22263477720409788   0.7931486716882185   0.5806693898091208   0.4014969138477898
0.9400350460179003   0.6886797418342318   0.9091003941026365   0.6058232649618833   0.9082370034159192   0.39441468820136394   0.4386717254627424   0.10009926316208069   0.5225090109530682   0.4372177726850274   0.4407328442861362   0.6322650335294709   0.8080204168003533   0.7609571801195326   0.6428968834652087   0.7005376014245287   0.07732981384594349   0.186747805694846   0.5830780466726703   0.9361428658109896   0.8546950366418457   0.39359913400662755   0.0024086568635496015   0.5346459519631999   0.9146599906239453   0.7049193921723957   0.09330826276091304   0.9288226870013165   0.006422987208026162   0.3105047039710318   0.6546365372981706   0.8287234238392359   0.48391397625495797   0.8732869312860044   0.21390369301203446   0.19645839030976497   0.6758935594546046   0.11232975116647179   0.5710068095468258   0.4959207888852363   0.5985637456086612   0.9255819454716258   0.9879287628741554   0.5597779230742466   0.7438687089668156   0.5319828114649983   0.9855201060106058   0.02513197111104675   0.8292087183428702   0.8270634192926024   0.8922118432496928   0.09630928410973016   0.8227857311348441   0.5165587153215706   0.23757530595152215   0.2675858602704943   0.3388717548798862   0.6432717840355662   0.023671612939487677   0.07112746996072931   0.6629781954252815   0.5309420328690944   0.4526648033926619   0.575206681075493
0.06441444981662035   0.6053600873974686   0.4647360405185064   0.015428758001246434   0.32054574084980475   0.07337727593247038   0.4792159345079006   0.9902967868901997   0.4913370225069345   0.24631385663986793   0.5870040912582077   0.8939875027804695   0.6685512913720904   0.7297551413182973   0.34942878530668564   0.6264016425099752   0.32967953649220416   0.08648335728273114   0.325757172367198   0.5552741725492459   0.6667013410669227   0.5555413244136368   0.873092368974536   0.9800674914737528   0.6022868912503023   0.9501812370161682   0.4083563284560296   0.9646387334725064   0.2817411504004975   0.8768039610836977   0.929140393948129   0.9743419465823068   0.7904041278935631   0.6304901044438298   0.34213630268992123   0.08035444380183725   0.12185283652147269   0.9007349631255325   0.9927075173832356   0.453952801291862   0.7921733000292686   0.8142516058428013   0.6669503450160377   0.8986786287426161   0.12547195896234584   0.2587102814291646   0.7938579760415015   0.9186111372688632   0.5231850677120435   0.30852904441299644   0.38550164758547195   0.9539724037963568   0.24144391731154596   0.4317250833292987   0.4563612536373429   0.9796304572140501   0.4510397894179829   0.8012349788854689   0.11422495094742169   0.8992760134122127   0.32918695289651023   0.9005000157599363   0.1215174335641861   0.44532321212035075
0.5370136528672417   0.08624840991713503   0.4545670885481485   0.5466445833777347   0.41154169390489587   0.8275381284879705   0.6607091125066469   0.6280334461088715   0.8883566261928524   0.519009084074974   0.2752074649211749   0.6740610423125146   0.6469127088813064   0.0872840007456753   0.8188462112838321   0.6944305850984647   0.1958729194633235   0.2860490218602064   0.7046212603364104   0.7951545716862518   0.8666859665668133   0.38554900610027004   0.5831038267722243   0.34983135956590106   0.32967231369957156   0.29930059618313504   0.12853673822407577   0.8031867761881664   0.9181306197946757   0.4717624676951646   0.46782762571742886   0.17515333007929496   0.029773993601823326   0.9527533836201906   0.19262016079625394   0.5010922877667803   0.38286128472051695   0.8654693828745154   0.3737739495124219   0.8066617026683157   0.18698836525719342   0.5794203610143088   0.6691526891760116   0.011507130982063823   0.32030239869038013   0.1938713549140388   0.08604886240378731   0.6616757714161627   0.9906300849908086   0.8945707587309037   0.9575121241797115   0.8584889952279964   0.07249946519613287   0.4228082910357392   0.4896844984622826   0.6833356651487014   0.04272547159430955   0.47005490741554856   0.29706433766602874   0.1822433773819211   0.6598641868737927   0.6045855245410333   0.9232903881536069   0.37558167471360543
0.4728758216165992   0.025165163526724404   0.2541376989775953   0.3640745437315416   0.15257342292621906   0.8312938086126855   0.16808883657380796   0.7023987723153788   0.1619433379354105   0.9367230498817818   0.21057671239409645   0.8439097770873825   0.08944387273927762   0.5139147588460427   0.7208922139318138   0.16057411193868112   0.04671840114496807   0.04385985143049403   0.42382787626578505   0.97833073455676   0.38685421427117545   0.4392743268894608   0.5005374881121782   0.6027490598431546   0.9139783926545763   0.41410916336273634   0.24639978913458294   0.23867451611161306   0.7614049697283571   0.5828153547500508   0.07831095256077497   0.5362757437962342   0.5994616317929466   0.646092304868269   0.8677342401666785   0.6923659667088518   0.5100177590536691   0.13217754602222634   0.14684202623486475   0.5317918547701705   0.463299357908701   0.08831769459173232   0.7230141499690796   0.5534611202134105   0.07644514363752557   0.6490433677022716   0.22247666185690146   0.9507120603702559   0.16246675098294933   0.2349342043395352   0.9760768727223185   0.7120375442586429   0.40106178125459213   0.6521188495894845   0.8977659201615436   0.17576180046240866   0.8016001494616455   0.0060265447212155205   0.03003167999486499   0.48339583375355694   0.29158239040797634   0.8738489986989891   0.8831896537600002   0.9516039789833863
0.8282830324992754   0.7855313041072569   0.16017550379092058   0.3981428587699758   0.7518378888617498   0.1364879364049853   0.9376988419340191   0.4474307983997199   0.5893711378788005   0.9015537320654501   0.9616219692117006   0.735393254141077   0.18830935662420833   0.24943488247596562   0.0638560490501571   0.5596314536786684   0.3867092071625629   0.2434083377547501   0.033824369055292104   0.0762356199251114   0.09512681675458654   0.36955933905576094   0.15063471529529185   0.12463164094172503   0.2668437842553112   0.5840280349485041   0.9904592115043713   0.7264887821717493   0.5150058953935613   0.4475400985435187   0.05276036957035217   0.27905798377202934   0.9256347575147609   0.5459863664780686   0.09113840035865155   0.5436647296309524   0.7373254008905525   0.296551484002103   0.02728235130849446   0.984033275952284   0.35061619372798963   0.05314314624735294   0.9934579822532024   0.9077976560271726   0.2554893769734031   0.6835838071915921   0.8428232669579105   0.7831660150854476   0.9886455927180919   0.09955577224308798   0.8523640554535392   0.05667723291369832   0.47363969732453054   0.6520156736995693   0.7996036858831871   0.777619249141669   0.5480049398097696   0.1060293072215006   0.7084652855245355   0.23395451951071664   0.8106795389192171   0.8094778232193975   0.681182934216041   0.24992124355843265
0.46006334519122744   0.7563346769720446   0.6877249519628387   0.34212358753126004   0.20457396821782436   0.07275086978045259   0.8449016850049281   0.5589575724458125   0.21592837549973243   0.9731950975373646   0.9925376295513889   0.5022803395321142   0.7422886781752018   0.32117942383779535   0.1929339436682019   0.7246610903904452   0.19428373836543222   0.21515011661629477   0.4844686581436664   0.4907065708797286   0.38360419944621515   0.4056722933968972   0.8032857239276254   0.24078532732129593   0.9235408542549877   0.6493376164248525   0.11556077196478669   0.8986617397900359   0.7189668860371633   0.5765867466444   0.2706590869598585   0.3397041673442234   0.5030385105374309   0.6033916491070354   0.27812145740846955   0.8374238278121092   0.760749832362229   0.28221222526924   0.08518751374026763   0.11276273742166404   0.5664660939967968   0.06706210865294526   0.6007188555966012   0.6220561665419355   0.18286189455058166   0.6613898152560481   0.7974331316689759   0.38127083922063953   0.25932104029559394   0.012052198831195496   0.6818723597041891   0.48260909943060365   0.5403541542584306   0.4354654521867955   0.4112132727443306   0.14290493208638025   0.037315643720999735   0.8320738030797601   0.1330918153358611   0.305481104274271   0.27656581135877073   0.5498615778105201   0.04790430159559346   0.192718366852607
0.710099717361974   0.4827994691575748   0.44718544599899224   0.5706622003106715   0.5272378228113923   0.8214096539015268   0.6497523143300165   0.189391361090032   0.2679167825157983   0.8093574550703313   0.9678799546258272   0.7067822616594284   0.7275626282573676   0.37389200288353575   0.5566666818814966   0.563877329573048   0.6902469845363679   0.5418181998037757   0.42357486654563553   0.25839622529877704   0.41368117317759723   0.9919566219932555   0.3756705649500421   0.06567785844617008   0.7035814558156233   0.5091571528356806   0.9284851189510498   0.4950156581354985   0.17634363300423103   0.6877474989341539   0.2787328046210334   0.30562429704546656   0.9084268504884327   0.8783900438638226   0.3108528499952061   0.5988420353860382   0.18086422223106505   0.5044980409802868   0.7541861681137095   0.034964705812990146   0.4906172376946971   0.9626798411765112   0.330611301568074   0.7765684805142131   0.07693606451709988   0.9707232191832557   0.9549407366180319   0.710890622068043   0.3733546087014766   0.461566066347575   0.026455617666982113   0.21587496393254446   0.19701097569724557   0.7738185674134211   0.7477228130459487   0.9102506668870779   0.2885841252088128   0.8954285235495985   0.43686996305074255   0.3114086315010397   0.1077199029777478   0.3909304825693117   0.682683794937033   0.27644392568804954
0.6171026652830507   0.42825064139280045   0.352072493368959   0.4998754451738365   0.5401666007659508   0.45752742220954473   0.3971317567509271   0.7889848231057934   0.16681199206447425   0.9959613558619697   0.370676139083945   0.573109859173249   0.9698010163672287   0.22214278844854857   0.6229533260379962   0.6628591922861711   0.6812168911584158   0.32671426489895006   0.18608336298725373   0.3514505607851314   0.573496988180668   0.9357837823296384   0.5033995680502207   0.07500663509708187   0.9563943228976173   0.507533140936838   0.15132707468126166   0.5751311899232454   0.4162277221316665   0.05000571872729326   0.7541953179303346   0.786146366817452   0.24941573006719225   0.05404436286532356   0.38351917884638953   0.213036507644203   0.27961471369996355   0.831901574416775   0.7605658528083933   0.5501773153580319   0.5983978225415477   0.505187309517825   0.5744824898211395   0.19872675457290054   0.024900834360879733   0.5694035271881865   0.07108292177091882   0.12372011947581865   0.06850651146326242   0.06187038625134855   0.9197558470896572   0.5485889295525732   0.6522787893315959   0.011864667524055295   0.16556052915932262   0.7624425627351212   0.4028630592644037   0.9578203046587317   0.7820413503129331   0.5494060550909182   0.12324834556444011   0.12591873024195674   0.021475497504539837   0.9992287397328863
0.5248505230228924   0.6207314207241318   0.44699300768340033   0.8005019851599857   0.4999496886620126   0.051327893535945274   0.3759100859124815   0.6767818656841671   0.4314431771987502   0.9894575072845967   0.45615423882282435   0.12819293613159388   0.7791643878671543   0.9775928397605415   0.2905937096635017   0.36575037339647265   0.3763013286027506   0.019772535101809693   0.5085523593505686   0.8163443183055544   0.2530529830383105   0.893853804859853   0.4870768618460288   0.8171155785726681   0.7282024600154181   0.27312238413572115   0.040083854162628454   0.01661359341268233   0.22825277135340546   0.22179449059977588   0.664173768250147   0.3398317277285152   0.7968095941546552   0.23233698331517916   0.20801952942732263   0.21163879159692134   0.017645206287500964   0.25474414355463776   0.9174258197638209   0.8458884182004487   0.6413438776847503   0.23497160845282805   0.4088734604132523   0.0295440998948943   0.3882908946464399   0.3411178035929751   0.9217965985672235   0.2124285213222262   0.6600884346310217   0.06799541945725393   0.8817127444045951   0.19581492790954386   0.4318356632776163   0.846200928857478   0.21753897615444812   0.8559832001810287   0.6350260691229611   0.6138639455422988   0.0095194467271255   0.6443444085841074   0.6173808628354601   0.35911980198766114   0.09209362696330457   0.7984559903836587
0.9760369851507097   0.12414819353483313   0.6832201665500522   0.7689118904887643   0.5877460905042698   0.783030389941858   0.7614235679828287   0.5564833691665381   0.9276576558732481   0.7150349704846041   0.8797108235782336   0.36066844125699427   0.49582199259563176   0.8688340416271261   0.6621718474237855   0.5046852410759656   0.8607959234726708   0.2549700960848272   0.65265240069666   0.8603408324918583   0.2434150606372106   0.895850294097166   0.5605587737333554   0.06188484210819967   0.2673780754865009   0.7717021005623329   0.8773386071833031   0.2929729516194354   0.679631984982231   0.9886717106204749   0.11591503920047445   0.7364895824528972   0.751974329108983   0.27363674013587075   0.2362042156222408   0.375821141195903   0.2561523365133512   0.4048026985087447   0.5740323681984553   0.8711359001199374   0.3953564130406805   0.14983260242391752   0.9213799675017953   0.010795067628079094   0.1519413524034699   0.2539823083267515   0.36082119376843985   0.9489102255198795   0.884563276916969   0.48228020776441866   0.48348258658513665   0.6559372739004441   0.204931291934738   0.4936084971439438   0.36756754738466224   0.9194476914475469   0.45295696282575504   0.21997175700807303   0.1313633317624214   0.5436265502516439   0.19680462631240384   0.8151690584993283   0.557330963563966   0.6724906501317065
0.8014482132717233   0.6653364560754108   0.6359509960621709   0.6616955825036274   0.6495068608682535   0.4113541477486593   0.27512980229373096   0.712785356983748   0.7649435839512845   0.9290739399842407   0.7916472157085943   0.0568480830833039   0.5600122920165465   0.43546544284029687   0.42407966832393207   0.13740039163575704   0.10705532919079139   0.21549368583222384   0.29271633656151064   0.5937738413841132   0.9102507028783875   0.4003246273328955   0.7353853729975446   0.9212831912524067   0.1088024896066642   0.7349881712574846   0.09943437693537373   0.2595876087487793   0.45929562873841073   0.32363402350882536   0.8243045746416428   0.5468022517650313   0.6943520447871263   0.39456008352458466   0.03265735893304848   0.48995416868172736   0.1343397527705799   0.9590946406842877   0.6085776906091164   0.35255377704597035   0.027284423579788518   0.7436009548520639   0.3158613540476058   0.7587799356618572   0.11703372070140097   0.3432763275191685   0.5804759810500613   0.8374967444094505   0.008231231094736776   0.6082881562616839   0.4810416041146875   0.5779091356606713   0.548935602356326   0.28465413275285845   0.6567370294730447   0.031106883895639963   0.8545835575691997   0.8900940492282738   0.6240796705399962   0.5411527152139126   0.7202438047986198   0.930999408543986   0.015501979930879822   0.18859893816794224
0.6929593812188313   0.18739845369192204   0.699640625883274   0.42981900250608507   0.5759256605174303   0.8441221261727536   0.11916464483321282   0.5923222580966345   0.5676944294226935   0.23583396991106978   0.6381230407185253   0.014413122435963283   0.018758827066367507   0.9511798371582113   0.9813860112454806   0.9833062385403233   0.16417526949716782   0.06108578792993752   0.35730634070548434   0.4421535233264107   0.443931464698548   0.13008637938595152   0.3418043607746045   0.2535545851584685   0.7509720834797168   0.9426879256940295   0.6421637348913305   0.8237355826523834   0.17504642296228642   0.09856579952127589   0.5229990900581176   0.23141332455574892   0.6073519935395929   0.8627318296102061   0.8848760493395923   0.21700020211978566   0.5885931664732253   0.9115519924519948   0.9034900380941118   0.23369396357946234   0.4244178969760576   0.8504662045220572   0.5461836973886274   0.7915404402530516   0.9804864322775095   0.7203798251361058   0.20437933661402283   0.5379858550945831   0.22951434879779284   0.7776918994420763   0.5622156017226924   0.7142502724421996   0.05446792583550642   0.6791260999208004   0.039216511664574696   0.48283694788645065   0.4471159322959135   0.8163942703105943   0.15434046232498236   0.265836745766665   0.8585227658226882   0.9048422778585995   0.2508504242308706   0.032142782187202686
0.4341048688466306   0.054376073336542194   0.7046667268422433   0.2406023419341511   0.45361843656912104   0.33399624820043644   0.5002873902282204   0.702616486839568   0.22410408777132818   0.5563043487583601   0.9380717885055281   0.9883662143973684   0.16963616193582176   0.8771782488375597   0.8988552768409533   0.5055292665109178   0.7225202296399083   0.06078397852696543   0.744514814515971   0.23969252074425274   0.8639974638172201   0.15594170066836593   0.49366439028510034   0.20754973855705006   0.42989259497058946   0.10156562733182375   0.7889976634428572   0.966947396622899   0.9762741584014685   0.7675693791313873   0.28871027321463666   0.2643309097833309   0.7521700706301403   0.21126503037302719   0.35063848470910863   0.2759646953859625   0.5825339086943185   0.33408678153546745   0.45178320786815523   0.7704354288750448   0.8600136790544103   0.273302803008502   0.7072683933521843   0.5307429081307921   0.9960162152371902   0.11736110234013608   0.21360400306708388   0.323193169573742   0.5661236202666007   0.015795475008312333   0.4246063396242268   0.35624577295084303   0.5898494618651323   0.248226095876925   0.1358960664095901   0.0919148631675121   0.837679391234992   0.03696106550389782   0.7852575817004814   0.8159501677815496   0.2551454825406735   0.7028742839684303   0.33347437383232625   0.04551473890650482
0.3951318034862632   0.4295714809599283   0.626205980480142   0.5147718307757128   0.399115588249073   0.31221037861979223   0.41260197741305815   0.1915786612019708   0.8329919679824722   0.2964149036114799   0.9879956377888314   0.8353328882511278   0.24314250611733998   0.04818880773455489   0.8520995713792413   0.7434180250836157   0.405463114882348   0.01122774223065707   0.06684198967875979   0.9274678573020662   0.1503176323416745   0.3083534582622267   0.7333676158464335   0.8819531183955612   0.7551858288554113   0.8787819773022985   0.10716163536629154   0.3671812876198485   0.3560702406063383   0.5665715986825062   0.6945596579532334   0.17560262641787766   0.5230782726238661   0.27015669507102624   0.706564020164402   0.3402697381667499   0.2799357665065261   0.22196788733647138   0.8544644487851608   0.5968517130831342   0.8744726516241781   0.21074014510581432   0.7876224591064009   0.6693838557810681   0.7241550192825036   0.9023866868435876   0.054254843259967434   0.7874307373855068   0.9689691904270923   0.02360470954128919   0.9470932078936759   0.4202494497656583   0.612898949820754   0.457033110858783   0.25253354994044247   0.24464682334778065   0.08982067719688794   0.18687641578775674   0.5459695297760404   0.9043770851810308   0.8098849106903618   0.9649085284512854   0.6915050809908796   0.30752537209789654
0.9354122590661837   0.7541683833454711   0.9038826218844787   0.6381415163168285   0.2112572397836802   0.8517816965018835   0.8496277786245112   0.8507107789313216   0.24228804935658788   0.8281769869605943   0.9025345707308353   0.4304613291656633   0.6293890995358339   0.37114387610181127   0.6500010207903929   0.1858145058178827   0.539568422338946   0.1842674603140545   0.10403149101435245   0.28143742063685195   0.7296835116485841   0.21935893186276914   0.4125264100234728   0.9739120485389554   0.7942712525824003   0.4651905485172981   0.5086437881389941   0.3357705322221269   0.5830140127987201   0.6134088520154146   0.6590160095144829   0.4850597532908052   0.34072596344213224   0.7852318650548203   0.7564814387836476   0.054598424125141876   0.7113368639062984   0.4140879889530091   0.10648041799325471   0.8687839183072592   0.17176844156735244   0.22982052863895455   0.0024489269789022645   0.5873464976704073   0.44208492991876835   0.010461596776185404   0.5899225169554294   0.6134344491314518   0.6478136773363681   0.5452710482588873   0.0812787288164353   0.277663916909325   0.06479966453764789   0.9318621962434728   0.42226271930195236   0.7926041636185198   0.7240737010955156   0.1466303311886524   0.6657812805183048   0.7380057394933779   0.01273683718921726   0.7325423422356434   0.5593008625250501   0.8692218211861187
0.8409683956218649   0.5027218135966888   0.5568519355461479   0.2818753235157115   0.3988834657030965   0.4922602168205034   0.9669294185907183   0.6684408743842596   0.7510697883667284   0.9469891685616161   0.8856506897742831   0.39077695747493457   0.6862701238290806   0.015126972318143347   0.46338797047233066   0.5981727938564149   0.962196422733565   0.868496641129491   0.7976066899540258   0.860167054363037   0.9494595855443476   0.13595429889384758   0.2383058274289758   0.9909452331769182   0.10849118992248283   0.6332324852971588   0.681453891882828   0.7090699096612068   0.7096077242193863   0.14097226847665537   0.7145244732921096   0.040629035276947174   0.9585379358526579   0.1939830999150393   0.8288737835178266   0.6498520778020126   0.2722678120235773   0.17885612759689595   0.3654858130454959   0.05167928394559775   0.3100713892900124   0.310359486467405   0.56787912309147   0.1915122295825608   0.3606118037456647   0.1744051875735574   0.3295732956624942   0.20056699640564257   0.2521206138231819   0.5411727022763987   0.6481194037796663   0.4914970867444358   0.5425128896037955   0.4002004337997433   0.9335949304875567   0.45086805146748865   0.5839749537511376   0.20621733388470398   0.10472114696973012   0.801015973665476   0.31170714172756037   0.027361206287808033   0.7392353339242342   0.7493366897198783
0.001635752437547948   0.7170017198204031   0.17135621083276426   0.5578244601373175   0.6410239486918832   0.5425965322468456   0.84178291517027   0.35725746373167494   0.3889033348687013   0.0014238299704469506   0.19366351139060378   0.8657603769872391   0.8463904452649058   0.6012233961707036   0.26006858090304713   0.41489232551975047   0.26241549151376814   0.3950060622859997   0.15534743393331701   0.6138763518542744   0.9507083497862078   0.36764485599819163   0.4161121000090828   0.864539662134396   0.9490725973486599   0.6506431361777887   0.24475588917631852   0.3067152019970786   0.3080486486567766   0.10804660393094302   0.4029729740060485   0.9494577382654037   0.9191453137880753   0.10662277396049608   0.20930946261544467   0.08369736127816456   0.0727548685231695   0.5053993777897924   0.9492408817123975   0.6688050357584141   0.8103393770094014   0.11039331550379272   0.7938934477790806   0.054928683904139707   0.8596310272231935   0.7427484595056011   0.3777813477699977   0.19038902176974362   0.9105584298745337   0.09210532332781243   0.13302545859367923   0.883673819772665   0.6025097812177571   0.9840587193968694   0.7300524845876307   0.9342160815072614   0.6833644674296818   0.8774359454363734   0.5207430219721861   0.8505187202290968   0.6106095989065123   0.37203656764658094   0.5715021402597885   0.18171368447068273
0.800270221897111   0.2616432521427882   0.7776086924807081   0.12678500056654302   0.9406391946739174   0.5188947926371872   0.3998273447107103   0.9363959787967994   0.03008076479938369   0.4267894693093747   0.2668018861170311   0.05272215902413434   0.4275709835816266   0.44273074991250533   0.5367494015294003   0.11850607751687295   0.7442065161519448   0.565294804476132   0.016006379557214213   0.2679873572877761   0.1335969172454325   0.19325823682955104   0.44450423929742566   0.08627367281709342   0.33332669534832154   0.9316149846867628   0.6668955468167176   0.9594886722505505   0.39268750067440417   0.4127201920495757   0.2670682021060073   0.02309269345375103   0.36260673587502046   0.985930722740201   0.00026631598897623016   0.9703705344296167   0.9350357522933939   0.5431999728276957   0.46351691445957593   0.8518644569127437   0.19082923614144903   0.9779051683515637   0.4475105349023617   0.5838770996249676   0.05723231889601654   0.7846469315220127   0.003006295604936056   0.49760342680787417   0.7239056235476949   0.8530319468352499   0.33611074878821845   0.5381147545573238   0.33121812287329083   0.44031175478567414   0.06904254668221114   0.5150220611035727   0.9686113869982704   0.45438103204547314   0.06877623069323492   0.544651526673956   0.033575634704876546   0.9111810592177775   0.605259316233659   0.6927870697612123
0.8427463985634275   0.9332758908662138   0.15774878133129727   0.1089099701362447   0.7855140796674109   0.1486289593442011   0.15474248572636123   0.6113065433283705   0.061608456119715965   0.29559701250895126   0.8186317369381427   0.07319178877104675   0.7303903332464251   0.8552852577232771   0.7495891902559316   0.558169727667474   0.7617789462481547   0.400904225677804   0.6808129595626967   0.013518200993517955   0.7282033115432782   0.4897231664600265   0.07555364332903772   0.3207311312323056   0.8854569129798506   0.5564472755938128   0.9178048619977405   0.21182116109606094   0.09994283331243971   0.4078183162496117   0.7630623762713792   0.6005146177676904   0.03833437719272375   0.1122213037406604   0.9444306393332365   0.5273228289966436   0.30794404394629865   0.2569360460173833   0.1948414490773048   0.9691531013291697   0.5461650976981439   0.8560318203395793   0.5140284895146081   0.9556349003356517   0.8179617861548657   0.3663086538795528   0.43847484618557037   0.6349037691033461   0.9325048731750151   0.80986137828574   0.52066998418783   0.42308260800728514   0.8325620398625754   0.4020430620361284   0.7576076079164508   0.8225679902395947   0.7942276626698516   0.28982175829546797   0.8131769685832143   0.295245161242951   0.48628361872355297   0.0328857122780847   0.6183355195059095   0.3260920599137814
0.940118521025409   0.1768538919385054   0.10430702999130141   0.3704571595781297   0.12215673487054332   0.8105452380589526   0.6658321838057311   0.7355533904747836   0.18965186169552825   0.0006838597732125812   0.1451621996179011   0.3124707824674985   0.3570898218329529   0.5986407977370842   0.3875545917014504   0.4899027922279038   0.5628621591631012   0.30881903944161626   0.574377623118236   0.19465763098495273   0.07657854043954829   0.2759333271635315   0.9560421036123266   0.8685655710711714   0.1364600194141392   0.09907943522502613   0.8517350736210252   0.49810841149304164   0.014303284543595907   0.28853419716607354   0.18590288981529413   0.762555021018258   0.8246514228480677   0.2878503373928609   0.040740690197393015   0.4500842385507596   0.4675616010151148   0.6892095396557767   0.6531860984959427   0.9601814463228557   0.9046994418520136   0.3803905002141605   0.07880847537770656   0.765523815337903   0.8281209014124652   0.10445717305062896   0.12276637176538   0.8969582442667318   0.691660881998326   0.005377737825602822   0.27103129814435484   0.39884983277369007   0.6773575974547301   0.7168435406595293   0.08512840832906071   0.636294811755432   0.8527061746066624   0.42899320326666834   0.044387718131667704   0.18621057320467246   0.38514457359154763   0.7397836636108917   0.3912016196357251   0.22602912688181667
0.4804451317395341   0.35939316339673116   0.3123931442580185   0.4605053115439136   0.6523242303270689   0.2549359903461022   0.1896267724926385   0.5635470672771818   0.9606633483287429   0.24955825252049937   0.9185954743482837   0.16469723450349183   0.2833057508740128   0.5327147118609701   0.8334670660192229   0.5284024227480598   0.43059957626735035   0.1037215085943017   0.7890793478875553   0.3421918495433873   0.045455002675802665   0.36393784498341003   0.3978777282518302   0.11616272266157067   0.5650098709362685   0.0045446815866789034   0.08548458399381169   0.6556574111176571   0.9126856406091997   0.7496086912405767   0.8958578115011732   0.09211034384047516   0.9520222922804568   0.5000504387200774   0.9772623371528895   0.9274131093369833   0.668716541406444   0.9673357268591073   0.14379527113366655   0.3990106865889235   0.23811696513909367   0.8636142182648056   0.3547159232461113   0.056818837045536176   0.192661962463291   0.4996763732813955   0.9568381949942811   0.9406561143839655   0.6276520915270225   0.4951316916947166   0.8713536110004694   0.28499870326630844   0.7149664509178228   0.7455230004541399   0.9754957994992962   0.1928883594258333   0.7629441586373661   0.24547256173406257   0.9982334623464068   0.26547525008885   0.0942276172309221   0.27813683487495533   0.8544381912127401   0.8664645634999264
0.8561106520918285   0.4145226166101498   0.49972226796662883   0.8096457264543903   0.6634486896285374   0.9148462433287543   0.5428840729723478   0.8689896120704248   0.03579659810151496   0.41971455163403765   0.6715304619718784   0.5839909088041163   0.3208301471836921   0.6741915511798978   0.6960346624725822   0.391102549378283   0.557885988546326   0.4287189894458352   0.6978012001261754   0.12562729928943303   0.46365837131540394   0.1505821545708799   0.8433630089134353   0.2591627357895066   0.6075477192235755   0.7360595379607301   0.3436407409468064   0.44951700933511635   0.9440990295950381   0.8212132946319759   0.8007566679744587   0.5805273972646916   0.9083024314935231   0.40149874299793825   0.1292262060025803   0.9965364884605753   0.587472284309831   0.7273071918180405   0.43319154352999817   0.6054339390822923   0.029586295763504956   0.2985882023722053   0.7353903434038228   0.47980663979285926   0.565927924448101   0.14800604780132537   0.8920273344903875   0.22064390400335268   0.9583802052245255   0.4119465098405952   0.5483865935435811   0.7711268946682364   0.014281175629487424   0.5907332152086193   0.7476299255691224   0.19059949740354476   0.10597874413596431   0.1892344722106811   0.618403719566542   0.1940630089429695   0.5185064598261333   0.46192728039264064   0.1852121760365439   0.5886290698606772
0.48892016406262834   0.16333907802043537   0.44982183263272113   0.10882243006781794   0.9229922396145274   0.015333030219109993   0.5577944981423336   0.8881785260644652   0.9646120343900019   0.6033865203785148   0.009407904598752537   0.11705163139622893   0.9503308587605144   0.012653305169895419   0.2617779790296301   0.9264521339926841   0.8443521146245501   0.8234188329592144   0.643374259463088   0.7323891250497147   0.3258456547984168   0.36149155256657367   0.4581620834265441   0.14376005518903745   0.8369254907357885   0.1981524745461383   0.008340250793822952   0.034937625121219514   0.9139332511212611   0.18281944432702832   0.45054575265148933   0.14675909905675424   0.9493212167312592   0.5794329239485135   0.4411378480527368   0.029707467660525316   0.9989903579707449   0.5667796187786182   0.1793598690231067   0.10325533366784116   0.15463824334619472   0.7433607858194038   0.5359856095600187   0.3708662086181265   0.8287925885477779   0.3818692332528301   0.0778235261334746   0.22710615342908905   0.9918670978119895   0.18371675870669182   0.06948327533965164   0.19216852830786954   0.07793384669072839   0.0008973143796635215   0.6189375226881623   0.045409429251115296   0.12861262995946915   0.42146439043114997   0.17779967463542554   0.01570196159058998   0.1296222719887243   0.8546847716525319   0.9984398056123188   0.9124466279227488
0.9749840286425296   0.11132398583312801   0.46245419605230015   0.5415804193046223   0.14619144009475168   0.7294547525802979   0.38463066991882555   0.31447426587553323   0.1543243422827622   0.545737993873606   0.31514739457917396   0.12230573756766372   0.07639049559203381   0.5448406794939425   0.6962098718910116   0.07689630831654842   0.9477778656325647   0.12337628906279254   0.5184101972555861   0.061194346725958436   0.8181555936438404   0.2686915174102607   0.5199703916432673   0.1487477188032096   0.8431715650013107   0.1573675315771327   0.057516195590967094   0.6071672994985873   0.696980124906559   0.42791277899683483   0.6728855256721415   0.29269303362305404   0.5426557826237969   0.8821747851232288   0.3577381310929676   0.17038729605539035   0.46626528703176306   0.3373341056292863   0.6615282592019559   0.09349098773884193   0.5184874213991983   0.21395781656649376   0.14311806194636983   0.03229664101288349   0.700331827755358   0.9452662991562331   0.6231476703031026   0.8835489222096738   0.8571602627540472   0.7878987675791004   0.5656314747121355   0.27638162271108657   0.1601801378474882   0.35998598858226555   0.8927459490399939   0.9836885890880325   0.6175243552236913   0.4778112034590367   0.5350078179470265   0.8133012930326421   0.15125906819192828   0.14047709782975043   0.8734795587450704   0.7198103052938002
0.6327716467927299   0.9265192812632567   0.7303614967987005   0.6875136642809168   0.9324398190373719   0.9812529821070236   0.107213826495598   0.8039647420712429   0.07527955628332468   0.19335421452792326   0.5415823517834625   0.5275831193601563   0.9150994184358365   0.8333682259456577   0.6488364027434685   0.5438945302721239   0.29757506321214516   0.355557022486621   0.11382858479644213   0.7305932372394817   0.1463159950202169   0.2150799246568706   0.24034902605137168   0.01078293194568147   0.513544348227487   0.2885606433936139   0.5099875292526711   0.3232692676647647   0.581104529190115   0.3073076612865903   0.4027737027570731   0.5193045255935219   0.5058249729067904   0.11395344675866706   0.8611913509736105   0.9917214062333656   0.5907255544709539   0.28058522081300935   0.21235494823014203   0.4478268759612417   0.2931504912588087   0.9250281983263883   0.09852636343369989   0.71723363872176   0.1468344962385918   0.7099482736695177   0.8581773373823282   0.7064507067760786   0.6332901480111048   0.42138763027590376   0.3481898081296571   0.38318143911131386   0.052185618820989786   0.11407996898931345   0.945416105372584   0.8638769135177919   0.5463606459141994   0.0001265222306463885   0.08422475439897348   0.8721555072844264   0.9556350914432455   0.7195413014176371   0.8718698061688315   0.42432863132318466
0.6624846001844369   0.7945131030912488   0.7733434427351316   0.7070949926014246   0.5156501039458451   0.08456482942173105   0.9151661053528034   0.0006442858253460258   0.8823599559347403   0.6631771991458273   0.5669762972231462   0.6174628467140322   0.8301743371137504   0.5490972301565138   0.6215601918505622   0.7535859331962402   0.283813691199551   0.5489707079258674   0.5373354374515887   0.8814304259118139   0.3281785997563055   0.8294294065082304   0.6654656312827573   0.45710179458862915   0.6656939995718686   0.03491630341698161   0.8921221885476257   0.7500068019872046   0.15004389562602358   0.9503514739952506   0.9769560831948224   0.7493625161618586   0.26768393969128335   0.2871742748494233   0.4099797859716761   0.13189966944782636   0.43750960257753296   0.7380770446929095   0.7884195941211138   0.37831373625158615   0.15369591137798194   0.18910633676704203   0.2510841566695251   0.4968833103397723   0.8255173116216765   0.35967693025881164   0.5856185253867678   0.03978151575114312   0.15982331204980785   0.32476062684183005   0.693496336839142   0.28977471376393854   0.009779416423784262   0.3744091528465795   0.7165402536443197   0.54041219760208   0.7420954767325009   0.0872348779971562   0.3065604676726436   0.40851252815425365   0.30458587415496796   0.3491578333042467   0.5181408735515297   0.030198791902667534
0.15088996277698602   0.16005149653720468   0.2670567168820046   0.5333154815628952   0.32537265115530956   0.800374566278393   0.6814381914952369   0.49353396581175213   0.1655493391055017   0.47561393943656294   0.9879418546560947   0.20375925204781356   0.15576992268171744   0.10120478658998348   0.271401601011775   0.6633470544457335   0.41367444594921654   0.013969908592827287   0.9648411333391315   0.2548345262914799   0.1090885717942486   0.6648120752885806   0.4467002597876017   0.22463573438881235   0.9581986090172626   0.5047605787513759   0.17964354290559706   0.6913202528259171   0.6328259578619531   0.7043860124729828   0.4982053514103602   0.197786287014165   0.4672766187564513   0.22877207303641992   0.5102634967542655   0.9940270349663515   0.31150669607473386   0.12756728644643642   0.23886189574249045   0.33067998052061787   0.8978322501255174   0.11359737785360914   0.274020762403359   0.07584545422913799   0.7887436783312687   0.4487853025650286   0.8273205026157573   0.8512097198403257   0.8305450693140062   0.9440247238136527   0.6476769597101603   0.1598894670144085   0.1977191114520531   0.23963871134066983   0.14947160829980005   0.9621031800002435   0.7304424926956018   0.010866638304249915   0.6392081115455346   0.968076145033892   0.4189357966208679   0.8832993518578135   0.40034621580304414   0.6373961645132742
0.5211035464953506   0.7697019740042044   0.12632545339968512   0.5615507102841362   0.7323598681640818   0.3209166714391758   0.2990049507839278   0.7103409904438105   0.9018147988500758   0.3768919476255231   0.6513279910737675   0.5504515234294021   0.7040956873980226   0.13725323628485328   0.5018563827739675   0.5883483434291585   0.9736531947024208   0.12638659798060337   0.8626482712284329   0.6202721983952665   0.554717398081553   0.24308724612278987   0.46230205542538877   0.9828760338819923   0.03361385158620241   0.4733852721185855   0.3359766020257037   0.42132532359785607   0.30125398342212056   0.15246860067940973   0.03697165124177587   0.7109843331540455   0.3994391845720448   0.7755766530538867   0.38564366016800833   0.1605328097246435   0.6953434971740222   0.6383234167690334   0.8837872773940408   0.572184466295485   0.7216903024716013   0.51193681878843   0.021139006165607953   0.9519122679002185   0.1669729043900483   0.2688495726656401   0.5588369507402192   0.9690362340182263   0.1333590528038459   0.7954643005470545   0.22286034871451552   0.5477109104203702   0.8321050693817253   0.6429956998676448   0.18588869747273964   0.8367265772663247   0.43266588480968055   0.8674190468137581   0.8002450373047313   0.6761937675416811   0.7373223876356584   0.22909563004472486   0.9164577599106905   0.10400930124619613
0.01563208516405706   0.7171588112562949   0.8953187537450825   0.15209703334597757   0.8486591807740087   0.44830923859065475   0.3364818030048633   0.18306079932775127   0.7153001279701628   0.6528449380436002   0.1136214542903478   0.6353498889073811   0.8831950585884375   0.009849238175955368   0.9277327568176081   0.7986233116410564   0.45052917377875695   0.14243019136219717   0.12748771951287688   0.12242954409937523   0.7132067861430986   0.9133345613174724   0.21102995960218646   0.018420242853179104   0.6975747009790415   0.19617575006117746   0.315711205857104   0.8663232095072015   0.8489155202050328   0.7478665114705226   0.9792294028522407   0.6832624101794503   0.13361539223486996   0.09502157342692248   0.8656079485618929   0.047912521272069235   0.25042033364643246   0.08517233525096711   0.9378751917442847   0.24928920963101286   0.7998911598676754   0.94274214388877   0.8103874722314078   0.12685966553163763   0.08668437372457687   0.029407582571297615   0.5993575126292214   0.10843942267845852   0.3891096727455353   0.8332318325101201   0.28364630677211744   0.24211621317125698   0.5401941525405025   0.08536532103959749   0.30441690391987675   0.5588538029918066   0.40657876030563256   0.990343747612675   0.43880895535798387   0.5109412817197375   0.15615842665920013   0.905171412361708   0.5009337636136991   0.2616520720887246
0.35626726679152465   0.962429268472938   0.6905462913822913   0.134792406557087   0.26958289306694777   0.9330216859016404   0.09118877875306988   0.026352983878628465   0.8804732203214124   0.09978985339152019   0.8075424719809524   0.7842367707073715   0.34027906778090994   0.014424532351922701   0.5031255680610758   0.2253829677155648   0.9337003074752773   0.0240807847392477   0.06431661270309187   0.7144416859958274   0.7775418808160772   0.1189093723775398   0.5633828490893927   0.4527896139071027   0.42127461402455263   0.15648010390460185   0.8728365577071014   0.31799720735001574   0.15169172095760483   0.2234584180029615   0.7816477789540316   0.29164422347138724   0.2712185006361924   0.12366856461144131   0.9741053069730792   0.5074074527640158   0.9309394328552825   0.10924403225951862   0.4709797389120034   0.28202448504845096   0.9972391253800051   0.08516324752027092   0.40666312620891154   0.5675827990526237   0.21969724456392786   0.9662538751427311   0.8432802771195188   0.11479318514552095   0.7984226305393752   0.8097737712381293   0.9704437194124174   0.7967959777955053   0.6467309095817704   0.5863153532351678   0.18879594045838574   0.505151754324118   0.375512408945578   0.46264678862372643   0.2146906334853066   0.9977443015601022   0.44457297609029556   0.35340275636420787   0.7437108945733032   0.7157198165116512
0.4473338507102904   0.26823950884393694   0.3370477683643917   0.14813701745902755   0.22763660614636258   0.3019856337012058   0.4937674912448729   0.0333438323135066   0.4292139756069873   0.4922118624630765   0.5233237718324556   0.23654785451800137   0.7824830660252169   0.9058965092279088   0.3345278313740699   0.7313961001938833   0.4069706570796389   0.44324972060418233   0.11983719788876326   0.7336517986337812   0.9623976809893434   0.08984696423997446   0.37612630331546004   0.017931982122129975   0.5150638302790529   0.8216074553960375   0.03907853495106837   0.8697949646631025   0.28742722413269034   0.5196218216948317   0.5453110437061954   0.8364511323495958   0.858213248525703   0.027409959231755182   0.021987271873739864   0.5999032778315945   0.0757301825004861   0.12151345000384642   0.68745944049967   0.868507177637711   0.6687595254208472   0.6782637293996641   0.5676222426109068   0.13485537900392985   0.7063618444315038   0.5884167651596897   0.19149593929544667   0.11692339688179988   0.1912980141524509   0.7668093097636521   0.1524174043443783   0.24712843221869746   0.9038707900197606   0.24718748806882038   0.6071063606381829   0.4106772998691016   0.045657541494057534   0.2197775288370652   0.585119088764443   0.8107740220375071   0.9699273589935714   0.09826407883321879   0.897659648264773   0.9422668443997961
0.30116783357272425   0.4200003494335547   0.33003740565386624   0.8074114653958663   0.5948059891412204   0.831583584273865   0.13854146635841957   0.6904880685140664   0.4035079749887695   0.06477427451021292   0.9861240620140412   0.44335963629536895   0.49963718496900894   0.8175867864413925   0.3790177013758584   0.03268233642626731   0.45397964347495146   0.5978092576043273   0.7938986126114154   0.22190831438876013   0.48405228448138   0.49954517877110854   0.8962389643466424   0.279641469988964   0.18288445090865574   0.07954482933755386   0.5662015586927761   0.4722300045930977   0.5880784617674354   0.24796124506368883   0.42766009233435653   0.7817419360790313   0.18457048677866583   0.1831869705534759   0.4415360303203153   0.33838229978366235   0.6849333018096568   0.36560018411208334   0.0625183289444569   0.305699963357395   0.23095365833470544   0.767790926507756   0.2686197163330415   0.0837916489686349   0.7469013738533254   0.2682457477366475   0.3723807519863991   0.8041501789796709   0.5640169229446697   0.18870091839909361   0.806179193293623   0.33192017438657323   0.9759384611772344   0.9407396733354048   0.3785191009592664   0.550178238307542   0.7913679743985685   0.7575527027819289   0.936983070638951   0.21179593852387957   0.10643467258891166   0.39195251866984554   0.8744647416944942   0.9060959751664845
0.8754810142542062   0.6241615921620896   0.6058450253614527   0.8223043261978497   0.1285796404008808   0.35591584442544205   0.2334642733750536   0.018154147218178734   0.5645627174562111   0.1672149260263484   0.4272850800814307   0.6862339728316055   0.5886242562789767   0.22647525269094362   0.04876597912216428   0.1360557345240636   0.7972562818804082   0.4689225499090147   0.11178290848321319   0.924259796000184   0.6908216092914966   0.0769700312391692   0.237318166788719   0.01816382083369946   0.8153405950372903   0.4528084390770797   0.6314731414272663   0.1958594946358498   0.6867609546364095   0.09689259465163767   0.3980088680522127   0.17770534741767108   0.12219823718019841   0.9296776686252892   0.9707237879707821   0.49147137458606555   0.5335739809012217   0.7032024159343456   0.9219578088486178   0.35541564006200194   0.7363176990208135   0.2342798660253309   0.8101749003654045   0.43115584406181795   0.04549608972931683   0.1573098347861617   0.5728567335766855   0.41299202322811845   0.2301554946920265   0.704501395709082   0.9413835921494192   0.21713252859226867   0.5433945400556169   0.6076088010574443   0.5433747240972066   0.03942718117459759   0.42119630287541854   0.6779311324321551   0.5726509361264245   0.547955806588532   0.8876223219741969   0.9747287164978095   0.6506931272778068   0.19254016652653008
0.1513046229533835   0.7404488504724785   0.8405182269124022   0.7613843224647121   0.10580853322406666   0.5831390156863168   0.2676614933357167   0.34839229923659365   0.8756530385320401   0.8786376199772348   0.32627790118629746   0.131259770644325   0.3322584984764232   0.27102881891979047   0.7829031770890909   0.0918325894697274   0.9110621956010047   0.5930976864876354   0.21025224096266637   0.5438767828811953   0.023439873626807745   0.6183689699898259   0.5595591136848596   0.3513366163546653   0.8721352506734242   0.8779201195173475   0.7190408867724574   0.5899522938899532   0.7663267174493575   0.2947811038310307   0.45137939343674066   0.24155999465335948   0.8906736789173174   0.41614348385379585   0.12510149225044323   0.11030022400903448   0.5584151804408942   0.14511466493400538   0.34219831516135235   0.018467634539307082   0.6473529848398896   0.55201697844637   0.13194607419868595   0.4745908516581117   0.6239131112130818   0.9336480084565439   0.5723869605138263   0.12325423530344644   0.7517778605396576   0.055727888939196536   0.853346073741369   0.5333019414134933   0.9854511430903   0.7609467851081659   0.40196668030462834   0.2917419467601338   0.09477746417298259   0.34480330125437003   0.2768651880541851   0.18144172275109935   0.5363622837320884   0.19968863632036465   0.9346668728928328   0.16297408821179227
0.8890092988921988   0.6476716578739947   0.8027207986941468   0.6883832365536805   0.26509618767911697   0.7140236494174507   0.2303338381803204   0.5651290012502341   0.5133183271394594   0.6582957604782541   0.37698776443895143   0.0318270598367408   0.5278671840491594   0.8973489753700883   0.9750210841343231   0.740085113076607   0.43308971987617684   0.5525456741157182   0.6981558960801381   0.5586433903255077   0.8967274361440885   0.3528570377953536   0.7634890231873053   0.39566930211371537   0.007718137251889643   0.7051853799213589   0.9607682244931585   0.7072860655600348   0.7426219495727726   0.9911617305039082   0.7304343863128381   0.14215706430980074   0.22930362243331326   0.33286597002565405   0.35344662187388665   0.11033000447305996   0.7014364383841538   0.4355169946555658   0.37842553773956356   0.370244891396453   0.26834671850797703   0.8829713205398475   0.6802696416594255   0.8116015010709453   0.3716192823638886   0.530114282744494   0.9167806184721202   0.41593219895722994   0.36390114511199895   0.824928902823135   0.9560123939789618   0.7086461333971951   0.6212791955392263   0.8337671723192268   0.2255780076661237   0.5664890690873944   0.391975573105913   0.5009012022935728   0.872131385792237   0.45615906461433436   0.6905391347217592   0.065384207638007   0.49370584805267353   0.08591417321788142
0.4221924162137821   0.18241288709815945   0.813436206393248   0.27431267214693605   0.050573133849893565   0.6522986043536655   0.8966555879211278   0.8583804731897061   0.6866719887378946   0.8273697015305304   0.940643193942166   0.14973433979251102   0.06539279319866836   0.9936025292113035   0.7150651862760423   0.5832452707051167   0.6734172200927553   0.4927013269177308   0.8429338004838053   0.1270862060907823   0.9828780853709962   0.42731711927972377   0.3492279524311317   0.04117203287290089   0.5606856691572141   0.24490423218156432   0.5357917460378837   0.7668593607259648   0.5101125353073205   0.5926056278278988   0.639136158116756   0.9084788875362587   0.8234405465694258   0.7652359262973685   0.69849296417459   0.7587445477437477   0.7580477533707575   0.7716333970860649   0.9834277778985476   0.17549927703863097   0.08463053327800213   0.27893207016833416   0.14049397741474243   0.04841307094784866   0.10175244790700597   0.8516149508886104   0.7912660249836108   0.007241038074947775   0.5410667787497919   0.6067107187070461   0.255474278945727   0.24038167734898297   0.03095424344247149   0.014105090879147226   0.6163381208289711   0.3319027898127243   0.20751369687304566   0.2488691645817788   0.9178451566543812   0.5731582420689766   0.4494659435022882   0.4772357674957139   0.9344173787558334   0.39765896503034565
0.36483541022428606   0.19830369732737976   0.7939234013410911   0.349245894082497   0.2630829623172801   0.3466887464387694   0.0026573763574803365   0.34200485600754926   0.7220161835674882   0.7399780277317233   0.7471830974117534   0.10162317865856627   0.6910619401250166   0.725872936852576   0.13084497658278227   0.7697203888458419   0.48354824325197104   0.4770037722707973   0.21299981992840117   0.19656214677686534   0.03408229974968281   0.9997680047750834   0.2785824411725677   0.7989031817465196   0.6692468895253967   0.8014643074477037   0.4846590398314766   0.4496572876640227   0.4061639272081166   0.45477556100893424   0.4820016634739963   0.10765243165647342   0.6841477436406285   0.714797533277211   0.7348185660622429   0.00602925299790716   0.9930858035156117   0.9889245964246348   0.6039735894794607   0.23630886415206517   0.5095375602636407   0.5119208241538376   0.39097376955105956   0.03974671737519983   0.4754552605139579   0.5121528193787541   0.11239132837849186   0.24084353562868016   0.8062083709885612   0.7106885119310505   0.6277322885470152   0.7911862479646575   0.40004444378044457   0.25591295092211624   0.1457306250730189   0.6835338163081841   0.7158967001398161   0.5411154176449053   0.41091205901077593   0.6775045633102769   0.7228108966242044   0.5521908212202704   0.8069384695313152   0.4411956991582117
0.21327333636056364   0.04026999706643288   0.41596469998025565   0.4014489817830119   0.7378180758466057   0.5281171776876787   0.3035733716017638   0.16060544615433175   0.9316097048580445   0.8174286657566282   0.6758410830547485   0.3694191981896743   0.5315652610775999   0.5615157148345119   0.5301104579817297   0.6858853818814902   0.8156685609377838   0.02040029718960665   0.11919839897095376   0.008380818571213294   0.09285766431357943   0.4682094759693362   0.31225992943963854   0.5671851194130015   0.8795843279530158   0.42793947890290335   0.8962952294593829   0.16573613762998968   0.14176625210641006   0.8998223012152246   0.5927218578576191   0.005130691475657933   0.21015654724836552   0.0823936354585964   0.9168807748028706   0.6357114932859836   0.6785912861707656   0.5208779206240844   0.3867703168211409   0.9498261114044935   0.8629227252329817   0.5004776234344778   0.26757191785018714   0.9414452928332802   0.7700650609194023   0.03226814746514159   0.9553119884105485   0.3742601734202786   0.8904807329663865   0.6043286685622382   0.059016758951165635   0.20852403579028894   0.7487144808599765   0.7045063673470137   0.4662949010935465   0.20339334431463102   0.538557933611611   0.6221127318884172   0.549414126290676   0.5676818510286473   0.8599666474408454   0.10123481126433281   0.16264380946953508   0.6178557396241539
0.9970439222078636   0.600757187829855   0.895071891619348   0.6764104467908737   0.22697886128846131   0.5684890403647134   0.9397599032087994   0.302150273370595   0.33649812832207476   0.9641603718024752   0.8807431442576338   0.09362623758030608   0.5877836474620983   0.2596540044554615   0.4144482431640873   0.8902328932656751   0.04922571385048738   0.6375412725670443   0.8650341168734114   0.32255104223702774   0.189259066409642   0.5363064613027114   0.7023903074038762   0.7046953026128739   0.19221514420177838   0.9355492734728564   0.8073184157845282   0.028284855822000247   0.9652362829133171   0.367060233108143   0.8675585125757288   0.7261345824514052   0.6287381545912423   0.40289986130566785   0.986815368318095   0.6325083448710991   0.040954507129143954   0.14324585685020635   0.5723671251540078   0.7422754516054241   0.9917287932786566   0.5057045842831621   0.7073330082805964   0.4197244093683963   0.8024697268690145   0.9693981229804506   0.0049427008767202055   0.7150291067555224   0.6102545826672362   0.0338488495075942   0.19762428509219196   0.6867442509335222   0.6450182997539191   0.6667886163994512   0.33006577251646313   0.9606096684821169   0.016280145162676868   0.26388875509378334   0.3432504041983681   0.3281013236110178   0.9753256380335329   0.12064289824357699   0.7708832790443604   0.5858258720055938
0.9835968447548763   0.6149383139604149   0.06355027076376392   0.16610146263719747   0.18112711788586178   0.6455401909799643   0.058607569887043715   0.45107235588167505   0.5708725352186256   0.61169134147237   0.8609832847948518   0.764328104948153   0.9258542354647065   0.9449027250729188   0.5309175122783886   0.8037184364660359   0.9095740903020295   0.6810139699791355   0.18766710808002052   0.4756171128550181   0.9342484522684966   0.5603710717355586   0.41678382903566014   0.8897912408494244   0.9506516075136203   0.9454327577751437   0.35323355827189623   0.7236897782122269   0.7695244896277585   0.2998925667951794   0.29462598838485254   0.27261742233055186   0.19865195440913297   0.6882012253228093   0.4336427035900008   0.5082893173823989   0.27279771894442656   0.7432985002498904   0.9027251913116121   0.704570880916363   0.363223628642397   0.06228453027075487   0.7150580832315916   0.22895376806134485   0.42897517637390037   0.5019134585351963   0.29827425419593145   0.3391625272119205   0.47832356886028005   0.5564807007600526   0.9450406959240353   0.6154727489996936   0.7087990792325215   0.2565881339648733   0.6504147075391827   0.34285532666914176   0.5101471248233885   0.568386908642064   0.21677200394918195   0.8345660092867428   0.237349405878962   0.8250884083921736   0.3140468126375698   0.12999512837037983
0.874125777236565   0.7628038781214187   0.5989887294059781   0.901041360309035   0.44515060086266467   0.2608904195862224   0.3007144752100467   0.5618788330971145   0.9668270320023846   0.7044097188261698   0.35567377928601146   0.9464060840974209   0.2580279527698631   0.4478215848612964   0.7052590717468288   0.6035507574282792   0.7478808279464746   0.8794346762192324   0.48848706779764683   0.7689847481415364   0.5105314220675126   0.05434626782705888   0.17444025516007705   0.6389896197711565   0.6364056448309475   0.29154238970564017   0.5754515257540989   0.7379482594621216   0.1912550439682829   0.030651970119417782   0.2747370505440522   0.1760694263650071   0.2244280119658983   0.3262422512932481   0.9190632712580407   0.22966334226758617   0.9664000591960352   0.8784206664319516   0.2138041995112119   0.626112584839307   0.21851923124956063   0.9989859902127192   0.725317131713565   0.8571278366977706   0.7079878091820481   0.9446397223856603   0.550876876553488   0.21813821692661398   0.07158216435110047   0.6530973326800201   0.9754253507993892   0.48018995746449233   0.8803271203828176   0.6224453625606023   0.700688300255337   0.3041205310994852   0.6558991084169192   0.29620311126735427   0.7816250289972964   0.07445718883189908   0.6894990492208841   0.41778244483540267   0.5678208294860845   0.44834460399259213
0.4709798179713235   0.4187964546226835   0.8425036977725193   0.5912167672948215   0.7629920087892754   0.47415673223702326   0.29162682121903133   0.3730785503682076   0.691409844438175   0.8210593995570031   0.3162014704196422   0.8928885929037153   0.8110827240553574   0.19861403699640087   0.6155131701643052   0.58876806180423   0.15518361563843813   0.9024109257290466   0.8338881411670088   0.5143108729723309   0.465684566417554   0.48462848089364396   0.26606731168092446   0.06596626897973878   0.9947047484462306   0.06583202627096048   0.4235636139084051   0.4747495016849172   0.23171273965695516   0.5916752940339373   0.1319367926893737   0.10167095131670963   0.5403028952187802   0.7706158944769341   0.8157353222697314   0.2087823584129944   0.7292201711634229   0.5720018574805332   0.2002221521054263   0.6200142966087644   0.5740365555249847   0.6695909317514865   0.36633401093841744   0.10570342363643348   0.10835198910743066   0.1849624508578426   0.10026669925749301   0.0397371546566947   0.11364724066120008   0.11913042458688212   0.676703085349088   0.5649876529717774   0.881934501004245   0.5274551305529449   0.5447662926597142   0.4633167016550679   0.34163160578546475   0.7568392360760108   0.7290309703899828   0.25453434324207347   0.612411434622042   0.18483737859547758   0.5288088182845565   0.6345200466333091
0.038374879097057224   0.515246446843991   0.16247480734613903   0.5288166229968756   0.9300228899896266   0.3302839959861484   0.06220810808864601   0.4890794683401809   0.8163756493284264   0.21115357139926627   0.38550502273955806   0.9240918153684035   0.9344411483241816   0.6836984408463214   0.8407387300798438   0.46077511371333557   0.5928095425387169   0.9268592047703106   0.11170775968986103   0.20624077047126207   0.9803981079166749   0.742021826174833   0.5828989414053046   0.571720723837953   0.9420232288196176   0.226775379330842   0.42042413405916557   0.04290410084107738   0.012000338829991122   0.8964913833446936   0.35821602597051955   0.5538246325008964   0.19562468950156464   0.6853378119454273   0.9727110032309615   0.6297328171324931   0.26118354117738307   0.0016393710991059584   0.13197227315111767   0.16895770341915747   0.6683739986386663   0.07478016632879537   0.02026451346125665   0.9627169329478954   0.6879758907219914   0.3327583401539624   0.43736557205595206   0.3909962091099424   0.7459526619023736   0.10598296082312036   0.01694143799678652   0.34809210826886505   0.7339523230723826   0.20949157747842675   0.658725412026267   0.7942674757679685   0.5383276335708179   0.5241537655329994   0.6860144087953055   0.1645346586354755   0.27714409239343485   0.5225143944338935   0.5540421356441878   0.9955769552163181
0.6087700937547685   0.44773422810509805   0.5337776221829311   0.03286002226842265   0.9207942030327773   0.11497588795113571   0.09641205012697909   0.6418638131584803   0.17484154113040354   0.008992927128015344   0.07947061213019257   0.29377170488961524   0.440889218058021   0.7995013496495886   0.4207452001039256   0.49950422912164666   0.902561584487203   0.27534758411658916   0.7347307913086201   0.33496957048617115   0.6254174920937683   0.7528331896826957   0.18068865566443226   0.3393926152698531   0.016647398338999704   0.30509896157759764   0.6469110334815011   0.3065325930014305   0.0958531953062225   0.19012307362646194   0.550498983354522   0.6646687798429503   0.921011654175819   0.1811301464984466   0.47102837122432945   0.370897074953335   0.480122436117798   0.38162879684885803   0.050283171120403834   0.8713928458316883   0.5775608516305949   0.10628121273226883   0.31555237981178375   0.5364232753455171   0.9521433595368266   0.35344802304957307   0.13486372414735145   0.19703066007566408   0.935495961197827   0.04834906147197543   0.48795269066585034   0.8904980670742336   0.8396427658916045   0.8582259878455135   0.9374537073113284   0.22582928723128343   0.9186311117157855   0.6770958413470669   0.46642533608699893   0.8549322122779484   0.4385086755979875   0.2954670444982089   0.4161421649665951   0.98353936644626
0.8609478239673926   0.18918583176594003   0.10058978515481136   0.44711609110074285   0.908804464430566   0.8357378087163669   0.9657260610074598   0.25008543102507874   0.9733085032327391   0.7873887472443916   0.47777337034160955   0.3595873639508451   0.13366573734113463   0.929162759398878   0.5403196630302811   0.13375807671956172   0.21503462562534917   0.25206691805181114   0.07389432694328224   0.2788258644416133   0.7765259500273617   0.9565998735536023   0.6577521619766872   0.2952864979953532   0.9155781260599691   0.7674140417876623   0.5571623768218757   0.8481704068946104   0.006773661629403097   0.9316762330712953   0.5914363158144159   0.5980849758695316   0.03346515839666404   0.14428748582690382   0.11366294547280638   0.2384976119186865   0.8997994210555293   0.21512472642802577   0.5733432824425252   0.10473953519912478   0.6847647954301802   0.9630578083762146   0.49944895549924295   0.8259136707575114   0.9082388454028185   0.006457934822612327   0.8416967935225559   0.5306271727621582   0.9926607193428495   0.23904389303495005   0.28453441670068   0.6824567658675479   0.9858870577134463   0.3073676599636547   0.6930981008862641   0.08437178999801621   0.9524218993167823   0.1630801741367509   0.5794351554134578   0.8458741780793297   0.05262247826125293   0.9479554477087251   0.006091872970932554   0.7411346428802049
0.36785768283107273   0.9848976393325105   0.5066429174716895   0.9152209721226935   0.45961883742825416   0.9784397045098981   0.6649461239491338   0.3845937993605353   0.4669581180854047   0.7393958114749482   0.3804117072484537   0.7021370334929874   0.48107106037195835   0.43202815151129337   0.6873136063621895   0.6177652434949712   0.528649161055176   0.26894797737454246   0.10787845094873176   0.7718910654156415   0.4760266827939231   0.3209925296658173   0.10178657797779922   0.030756422535436544   0.10816899996285036   0.3360948903333068   0.5951436605061097   0.11553545041274306   0.6485501625345962   0.3576551858234086   0.9301975365569759   0.7309416510522078   0.1815920444491915   0.6182593743484605   0.5497858293085223   0.02880461755922039   0.7005209840772332   0.18623122283716712   0.8624722229463326   0.4110393740642492   0.1718718230220572   0.9172832454626246   0.7545937719976009   0.6391483086486077   0.6958451402281342   0.5962907157968073   0.6528071940198017   0.6083918861131712   0.5876761402652838   0.2601958254635005   0.057663533513692064   0.4928564357004281   0.9391259777306875   0.9025406396400919   0.12746599695671615   0.7619147846482203   0.7575339332814961   0.2842812652916314   0.577680167648194   0.7331101670889999   0.05701294920426287   0.09805004245446426   0.7152079447018612   0.3220707930247507
0.8851411261822056   0.18076679699183962   0.9606141727042603   0.682922484376143   0.18929598595407154   0.5844760811950324   0.30780697868445867   0.07453059826297186   0.6016198456887878   0.3242802557315318   0.2501434451707666   0.5816741625625438   0.6624938679581003   0.42173961609143995   0.12267744821405042   0.8197593779143235   0.9049599346766042   0.1374583507998086   0.5449972805658565   0.08664921082532362   0.8479469854723413   0.03940830834534433   0.8297893358639952   0.7645784178005729   0.9628058592901356   0.8586415113535047   0.8691751631597349   0.08165593342442991   0.773509873336064   0.2741654301584724   0.5613681844752763   0.0071253351614580475   0.1718900276472763   0.9498851744269405   0.31122473930450967   0.4254511725989143   0.5093961596891761   0.5281455583355006   0.18854729109045923   0.6056917946845908   0.6044362250125719   0.390687207535692   0.6435500105246027   0.5190425838592672   0.7564892395402306   0.3512788991903477   0.8137606746606075   0.7544641660586943   0.793683380250095   0.49263738783684297   0.9445855115008727   0.6728082326342644   0.020173506914030866   0.2184719576783706   0.3832173270255964   0.6656828974728063   0.8482834792667546   0.26858678325143004   0.07199258772108678   0.240231724873892   0.3388873195775785   0.7404412249159293   0.8834452966306275   0.6345399301893012
0.7344510945650067   0.34975401738023737   0.23989528610602484   0.11549734633003408   0.9779618550247761   0.9984751181898897   0.4261346114454173   0.36103318027133985   0.18427847477468112   0.5058377303530467   0.48154909994454465   0.6882249476370755   0.16410496786065024   0.28736577267467606   0.09833177291894822   0.02254205016426925   0.3158214885938957   0.01877898942324606   0.026339185197861437   0.7823103252903773   0.9769341690163171   0.2783377645073167   0.14289388856723387   0.147770395101076   0.2424830744513105   0.9285837471270793   0.902998602461209   0.032273048771041916   0.26452121942653445   0.9301086289371896   0.47686399101579174   0.6712398684997021   0.08024274465185334   0.42427089858414296   0.995314891071247   0.9830149208626265   0.9161377767912031   0.13690512590946688   0.8969831181522988   0.9604728706983573   0.6003162881973074   0.11812613648622083   0.8706439329544374   0.17816254540798004   0.6233821191809903   0.8397883719789042   0.7277500443872036   0.030392150306904047   0.3808990447296798   0.9112046248518249   0.8247514419259945   0.9981191015358621   0.1163778253031453   0.9810959959146353   0.3478874509102028   0.32687923303616007   0.03613508065129196   0.5568250973304922   0.3525725598389557   0.3438643121735335   0.11999730386008886   0.4199199714210254   0.4555894416866569   0.38339144147517623
0.5196810156627815   0.30179383493480455   0.5849455087322195   0.2052288960671962   0.8962988964817912   0.46200546295590034   0.8571954643450159   0.17483674576029215   0.5153998517521114   0.5508008381040755   0.03244402241902144   0.17671764422443   0.3990220264489661   0.5697048421894403   0.6845565715088187   0.84983841118827   0.36288694579767417   0.012879744858948022   0.33198401166986297   0.5059740990147364   0.24288964193758528   0.5929597734379226   0.8763945699832061   0.12258265753956017   0.7232086262748039   0.2911659385031181   0.2914490612509866   0.917353761472364   0.8269097297930127   0.8291604755472177   0.43425359690597065   0.7425170157120718   0.3115098780409013   0.2783596374431423   0.4018095744869492   0.5657993714876418   0.9124878515919351   0.708654795253702   0.7172530029781305   0.7159609602993718   0.549600905794261   0.695775050394754   0.3852689913082676   0.20998686128463545   0.30671126385667574   0.1028152769568313   0.5088744213250616   0.08740420374507528   0.5835026375818719   0.8116493384537132   0.21742536007407495   0.1700504422727113   0.7565929077888592   0.9824888629064954   0.7831717631681043   0.4275334265606395   0.44508302974795794   0.7041292254633531   0.3813621886811551   0.8617340550729976   0.5325951781560228   0.9954744302096511   0.6641091857030246   0.14577309477362577
0.9829942723617617   0.29969937981489714   0.27884019439475694   0.9357862334889904   0.676283008505086   0.19688410285806585   0.7699657730696954   0.8483820297439151   0.0927803709232141   0.38523476440435267   0.5525404129956205   0.6783315874712037   0.3361874631343549   0.4027459014978573   0.7693686498275162   0.2507981609105643   0.891104433386397   0.6986166760345042   0.38800646114636106   0.3890641058375666   0.35850925523037425   0.703142245824853   0.7238972754433365   0.24329101106394085   0.3755149828686125   0.4034428660099558   0.4450570810485795   0.30750477757495054   0.6992319743635265   0.20655876315188998   0.6750913079788841   0.4591227478310355   0.6064516034403123   0.8213239987475374   0.12255089498326363   0.7807911603598318   0.27026414030595747   0.41857809724968004   0.3531822451557475   0.5299929994492675   0.37915970691956047   0.7199614212151759   0.9651757840093864   0.14092889361170086   0.020650451689186274   0.01681917539032292   0.24127850856604993   0.89763788254776   0.6451354688205738   0.6133763093803671   0.7962214275174704   0.5901331049728095   0.9459034944570474   0.4068175462284771   0.12113011953858632   0.13101035714177395   0.3394518910167349   0.5854935474809397   0.9985792245553227   0.3502191967819422   0.06918775071077746   0.16691545023125975   0.6453969793995752   0.8202261973326747
0.690028043791217   0.44695402901608383   0.6802211953901888   0.6792973037209739   0.6693775921020307   0.4301348536257609   0.43894268682413884   0.7816594211732139   0.024242123281456897   0.8167585442453938   0.6427212593066685   0.19152631620040436   0.0783386288244096   0.40994099801691675   0.5215911397680821   0.060515959058630414   0.7388867378076747   0.8244474505359769   0.5230119152127594   0.7102967622766883   0.6696989870968972   0.6575320003047171   0.8776149358131842   0.8900705649440136   0.9796709433056803   0.21057797128863337   0.19739374042299537   0.21077326122303977   0.3102933512036496   0.7804431176628724   0.7584510535988566   0.42911384004982595   0.2860512279221927   0.9636845734174786   0.1157297942921881   0.2375875238494216   0.20771259909778308   0.553743575400562   0.594138654524106   0.1770715647907912   0.4688258612901084   0.729296124864585   0.0711267393113466   0.46677480251410297   0.7991268741932112   0.07176412455986779   0.1935118034981624   0.5767042375700894   0.8194559308875309   0.8611861532712344   0.996118063075167   0.3659309763470496   0.5091625796838813   0.08074303560836195   0.2376670094763105   0.9368171362972236   0.22311135176168867   0.11705846219088331   0.12193721518412241   0.699229612447802   0.015398752663905588   0.5633148867903214   0.5277985606600164   0.5221580476570108
0.5465728913737972   0.8340187619257364   0.4566718213486698   0.05538324514290786   0.747446017180586   0.7622546373658686   0.2631600178505074   0.4786790075728185   0.9279900862930551   0.9010684840946342   0.2670419547753403   0.11274803122576892   0.4188275066091737   0.8203254484862723   0.02937494529902983   0.1759308949285453   0.19571615484748506   0.703266986295389   0.9074377301149075   0.4767012824807433   0.18031740218357947   0.13995209950506757   0.379639169454891   0.9545432348237325   0.6337445108097823   0.3059333375793311   0.9229673481062212   0.8991599896808247   0.8862984936291963   0.5436787002134625   0.6598073302557138   0.42048098210800616   0.9583084073361412   0.6426102161188283   0.3927653754803735   0.30773295088223723   0.5394809007269675   0.822284767632556   0.36339043018134365   0.13180205595369193   0.3437647458794824   0.11901778133716703   0.45595270006643623   0.6551007734729486   0.16344734369590294   0.9790656818320995   0.07631353061154521   0.7005575386492161   0.5297028328861206   0.6731323442527684   0.153346182505324   0.8013975489683915   0.6434043392569243   0.12945364403930587   0.4935388522496102   0.3809165668603854   0.6850959319207831   0.4868434279204776   0.10077347676923672   0.07318361597814815   0.14561503119381566   0.6645586602879217   0.7373830465878931   0.9413815600244562
0.8018502853143332   0.5455408789507545   0.2814303465214569   0.28628078655150757   0.6384029416184303   0.5664751971186551   0.20511681590991165   0.5857232479022915   0.10870010873230965   0.8933428528658868   0.05177063340458764   0.7843256989338999   0.4652957694753853   0.7638892088265808   0.5582317811549774   0.40340913207351453   0.7801998375546022   0.2770457809061033   0.45745830438574075   0.3302255160953664   0.6345848063607865   0.6124871206181817   0.7200752577978476   0.38884395607091016   0.8327345210464533   0.06694624166742712   0.43864491127639077   0.1025631695194026   0.19433157942802298   0.500471044548772   0.23352809536647914   0.5168399216171111   0.08563147069571332   0.6071281916828852   0.18175746196189152   0.7325142226832112   0.620335701220328   0.8432389828563044   0.6235256808069141   0.32910509060969667   0.8401358636657259   0.5661932019502011   0.16606737642117333   0.9988795745143303   0.2055510573049394   0.9537060813320194   0.44599211862332566   0.6100356184434201   0.3728165362584861   0.8867598396645923   0.007347207346934884   0.5074724489240175   0.17848495683046314   0.38628879511582026   0.7738191119804557   0.9906325273069063   0.09285348613474982   0.779160603432935   0.5920616500185643   0.2581183046236951   0.4725177849144218   0.9359216205766306   0.9685359692116502   0.9290132140139984
0.6323819212486959   0.3697284186264296   0.8024685927904769   0.9301336394996682   0.4268308639437565   0.41602233729441024   0.35647647416715117   0.32009802105624807   0.05401432768527042   0.5292624976298179   0.3491292668202163   0.8126255721322305   0.8755293708548073   0.14297370251399774   0.5753101548397606   0.8219930448253242   0.7826758847200574   0.36381309908106274   0.9832485048211963   0.5638747402016291   0.3101580998056357   0.4278914785044321   0.014712535609546142   0.6348615261876307   0.6777761785569397   0.05816305987800253   0.2122439428190693   0.7047278866879625   0.2509453146131832   0.6421407225835923   0.8557674686519181   0.3846298656317144   0.1969309869279128   0.11287822495377434   0.5066382018317018   0.5720042934994839   0.3214016160731055   0.9699045224397767   0.9313280469919413   0.7500112486741597   0.538725731353048   0.6060914233587139   0.948079542170745   0.18613650847253055   0.2285676315474124   0.17819994485428176   0.9333670065611989   0.5512749822848999   0.5507914529904726   0.12003688497627922   0.7211230637421295   0.8465470955969374   0.2998461383772894   0.4778961623926869   0.8653555950902114   0.46191722996522294   0.1029151514493766   0.3650179374389126   0.35871739325850954   0.8899129364657391   0.7815135353762711   0.395113414999136   0.42738934626656827   0.1399016877915794
0.242787804023223   0.7890219916404221   0.47930980409582324   0.9537651793190489   0.014220172475810608   0.6108220467861404   0.5459427975346244   0.40249019703414896   0.463428719485338   0.49078516180986115   0.8248197337924948   0.5559431014372116   0.16358258110804855   0.012888999417174241   0.9594641387022834   0.09402587147198864   0.06066742965867195   0.6478710619782617   0.6007467454437738   0.20411293500624958   0.2791538942824009   0.25275764697912567   0.17335739917720555   0.06421124721467014   0.03636609025917786   0.4637356553387036   0.6940475950813824   0.11044606789562128   0.022145917783367258   0.8529136085525632   0.14810479754675795   0.7079558708614723   0.5587171982980292   0.36212844674270206   0.3232850637542632   0.1520127694242607   0.3951346171899807   0.3492394473255278   0.3638209250519798   0.05798689795227206   0.3344671875313088   0.7013683853472662   0.763074179608206   0.8538739629460225   0.055313293248907915   0.44861073836814047   0.5897167804310004   0.7896627157313524   0.018947202989730048   0.9848750830294369   0.8956691853496181   0.6792166478357311   0.9968012852063628   0.13196147447687367   0.7475643878028602   0.9712607769742587   0.4380840869083335   0.7698330277341716   0.424279324048597   0.819248007549998   0.04294946971835277   0.4205935804086438   0.06045839899661718   0.761261109597726
0.708482282187044   0.7192251950613777   0.2973842193884112   0.9073871466517035   0.653168988938136   0.2706144566932372   0.7076674389574107   0.11772443092035115   0.6342217859484061   0.2857393736638003   0.8119982536077927   0.4385077830846201   0.6374205007420433   0.15377789918692664   0.06443386580493247   0.4672470061103613   0.19933641383370973   0.383944871452755   0.6401545417563355   0.6479989985603632   0.15638694411535697   0.9633512910441112   0.5796961427597183   0.8867378889626373   0.44790466192831296   0.24412609598273352   0.2823119233713071   0.9793507423109338   0.7947356729901769   0.9735116392894964   0.5746444844138964   0.8616263113905827   0.1605138870417709   0.687772265625696   0.7626462308061037   0.4231185283059625   0.5230933862997277   0.5339943664387693   0.6982123650011712   0.9558715221956012   0.3237569724660179   0.15004949498601433   0.058057823244835785   0.307872523635238   0.16737002835066095   0.18669820394190312   0.47836168048511746   0.4211346346726007   0.7194653664223479   0.9425721079591696   0.19604975711381037   0.44178389236166693   0.924729693432171   0.9690604686696732   0.621405272699914   0.5801575809710843   0.7642158063904002   0.2812882030439773   0.8587590418938102   0.15703905266512175   0.2411224200906725   0.7472938366052079   0.16054667689263896   0.20116753046952052
0.9173654476246546   0.5972443416191936   0.10248885364780318   0.8932950068342825   0.7499954192739936   0.4105461376772905   0.6241271731626857   0.47216037216168183   0.03053005285164568   0.46797402971812085   0.42807741604887534   0.030376479800014927   0.10580035941947463   0.4989135610484476   0.8066721433489613   0.4502188988289306   0.3415845530290745   0.21762535800447033   0.9479131014551512   0.2931798461638089   0.10046213293840196   0.47033152139926243   0.7873664245625122   0.09201231569428839   0.18309668531374737   0.8730871797800688   0.684877570914709   0.19871730886000585   0.43310126603975374   0.46254104210277835   0.0607503977520233   0.726556936698324   0.40257121318810807   0.9945670123846575   0.632672981703148   0.6961804568983091   0.29677085376863344   0.49565345133620986   0.8260008383541866   0.24596155806937844   0.9551863007395589   0.27802809333173956   0.8780877368990355   0.9527817119055696   0.854724167801157   0.8076965719324771   0.09072131233652331   0.8607693962112811   0.6716274824874097   0.9346093921524083   0.40584374142181434   0.6620520873512753   0.2385262164476559   0.47206835004962994   0.345093343669791   0.9354951506529513   0.8359550032595479   0.4775013376649725   0.712420361966643   0.23931469375464223   0.5391841494909144   0.9818478863287626   0.8864195236124565   0.9933531356852637
0.5839978487513554   0.7038197929970231   0.008331786713420955   0.04057142377969424   0.7292736809501985   0.896123221064546   0.9176104743768977   0.1798020275684131   0.057646198462788845   0.9615138289121377   0.5117667329550833   0.5177499402171378   0.8191199820151329   0.4894454788625077   0.16667338928529232   0.5822547895641865   0.9831649787555852   0.011944141197535242   0.45425302731864925   0.34294009580954427   0.4439808292646707   0.030096254868772633   0.5678335037061928   0.3495869601242805   0.8599829805133152   0.3262764618717496   0.5595017169927718   0.30901553634458623   0.1307092995631168   0.4301532408072036   0.6418912426158743   0.12921350877617316   0.07306310110032796   0.4686394118950659   0.13012450966079092   0.6114635685590354   0.253943119085195   0.9791939330325582   0.9634511203754986   0.02920877899484889   0.27077814032960984   0.967249791835023   0.5091980930568494   0.6862686831853047   0.8267973110649391   0.9371535369662504   0.9413645893506565   0.3366817230610241   0.9668143305516239   0.6108770750945007   0.38186287235788463   0.0276661867164379   0.8361050309885071   0.18072383428729719   0.7399716297420104   0.8984526779402647   0.7630419298881791   0.7120844223922312   0.6098471200812194   0.28698910938122935   0.5090988108029841   0.732890489359673   0.6463959997057208   0.2577803303863805
0.23832067047337427   0.76564069752465   0.13719790664887155   0.5715116472010758   0.4115233594084351   0.8284871605583998   0.19583331729821507   0.23482992414005172   0.44470902885681124   0.21761008546389896   0.8139704449403304   0.20716373742361383   0.6086039978683042   0.03688625117660176   0.07399881519832008   0.3087110594833491   0.845562067980125   0.3248018287843705   0.46415169511710064   0.0217219501021197   0.33646325717714093   0.5919113394246974   0.8177556954113797   0.7639416197157393   0.09814258670376665   0.8262706419000474   0.6805577887625082   0.19242997251466337   0.6866192272953315   0.9977834813416476   0.48472447146429315   0.9576000483746117   0.2419101984385203   0.7801733958777487   0.6707540265239627   0.7504363109509978   0.6333062005702161   0.743287144701147   0.5967552113256426   0.44172525146764874   0.7877441325900911   0.4184853159167764   0.132603516208542   0.42000330136552905   0.4512808754129502   0.826573976492079   0.3148478207971622   0.6560616816497898   0.3531382887091835   0.00030333459203159643   0.6342900320346541   0.46363170913512647   0.666519061413852   0.002519853250383953   0.1495655605703609   0.5060316607605149   0.4246088629753317   0.22234645737263525   0.4788115340463982   0.755595349809517   0.7913026624051156   0.4790593126714883   0.8820563227207556   0.31387009834186824
0.003558529815024485   0.0605739967547119   0.7494528065122136   0.8938667969763392   0.5522776544020743   0.23400002026263292   0.43460498571505135   0.23780511532654933   0.19913936569289079   0.23369668567060134   0.8003149536803973   0.7741734061914228   0.5326203042790388   0.2311768324202174   0.6507493931100364   0.268141745430908   0.1080114413037071   0.008830375047582117   0.17193785906363818   0.512546395621391   0.3167087788985915   0.5297710623760938   0.28988153634288255   0.19867629727952277   0.31315024908356703   0.46919706562138186   0.5404287298306689   0.3048095003031836   0.7608725946814927   0.23519704535874894   0.10582374411561762   0.06700438497663425   0.5617332289886019   0.0015003596881476198   0.30550879043522033   0.29283097878521136   0.029112924709563143   0.7703235272679303   0.654759397325184   0.024689233354303366   0.9211014834058561   0.7614931522203481   0.4828215382615458   0.5121428377329124   0.6043927045072646   0.23172208984425435   0.1929400019186632   0.31346654045338956   0.2912424554236975   0.7625250242228725   0.6525112720879942   0.00865704015020601   0.5303698607422047   0.5273279788641235   0.5466875279723766   0.9416526551735718   0.9686366317536028   0.5258276191759759   0.24117873753715627   0.6488216763883604   0.9395237070440396   0.7555040919080457   0.5864193402119723   0.624132443034057
0.018422223638183622   0.9940109396876975   0.10359780195042657   0.11198960530114467   0.4140295191309191   0.7622888498434431   0.9106578000317633   0.798523064847755   0.12278706370722163   0.9997638256205708   0.25814652794376913   0.7898660246975491   0.5924172029650169   0.47243584675644723   0.7114589999713926   0.8482133695239773   0.6237805712114141   0.9466082275804714   0.47028026243423626   0.19939169313561692   0.6842568641673744   0.19110413567242568   0.883860922222264   0.5752592501015599   0.6658346405291908   0.19709319598472813   0.7802631202718374   0.4632696448004152   0.25180512139827166   0.43480434614128494   0.869605320240074   0.6647465799526602   0.12901805769105004   0.43504052052071424   0.6114587922963048   0.8748805552551111   0.5366008547260331   0.9626046737642671   0.8999997923249122   0.026667185731133778   0.9128202835146191   0.01599644618379572   0.42971952989067597   0.8272754925955169   0.2285634193472447   0.82489231051137   0.545858607668412   0.252016242493957   0.5627287788180539   0.6277991145266419   0.7655954873965747   0.7887465976935417   0.31092365741978223   0.19299476838535695   0.8959901671565007   0.12400001774088162   0.1819055997287322   0.7579542478646427   0.2845313748601958   0.24911946248577055   0.6453047450026991   0.7953495741003757   0.3845315825352835   0.22245227675463677
0.7324844614880799   0.77935312791658   0.9548120526446076   0.3951767841591199   0.5039210421408352   0.9544608174052099   0.4089534449761955   0.14316054166516293   0.9411922633227813   0.326661702878568   0.6433579575796209   0.3544139439716211   0.630268605902999   0.13366693449321104   0.7473677904231202   0.23041392623073953   0.4483630061742669   0.3757126866285683   0.4628364155629244   0.981294463744969   0.8030582611715679   0.5803631125281926   0.07830483302764085   0.7588421869903322   0.07057379968348794   0.8010099846116127   0.12349278038303332   0.3636654028312123   0.5666527575426528   0.8465491672064028   0.7145393354068378   0.22050486116604937   0.6254604942198714   0.5198874643278348   0.071181377827217   0.8660909171944282   0.9951918883168723   0.38622052983462374   0.3238135874040968   0.6356769909636887   0.5468288821426055   0.010507843206055424   0.8609771718411724   0.6543825272187197   0.7437706209710376   0.4301447306778628   0.7826723388135316   0.8955403402283876   0.6731968212875497   0.6291347460662501   0.6591795584304982   0.5318749373971753   0.10654406374489693   0.7825855788598473   0.9446402230236605   0.3113700762311259   0.4810835695250255   0.26269811453201247   0.8734588451964435   0.4452791590366976   0.4858916812081532   0.8764775846973888   0.5496452577923466   0.809602168073009
0.9390627990655478   0.8659697414913333   0.6886680859511741   0.15521964085428921   0.19529217809451016   0.4358250108134705   0.9059957471376426   0.25967930062590167   0.5220953568069605   0.8066902647472205   0.24681618870714434   0.7278043632287264   0.41555129306206356   0.024104685887373183   0.30217596568348387   0.4164342869976006   0.934467723537038   0.7614065713553607   0.42871712048704047   0.971155127960903   0.44857604232888487   0.8849289866579719   0.8790718626946938   0.16155295988789398   0.5095132432633371   0.018959245166638647   0.1904037767435197   0.00633331903360476   0.3142210651688269   0.5831342343531681   0.2844080296058771   0.7466540184077031   0.7921257083618664   0.7764439696059476   0.03759184089873276   0.018849655178976632   0.3765744152998028   0.7523392837185745   0.7354158752152489   0.6024153681813761   0.44210669176276474   0.9909327123632138   0.3066987547282084   0.6312602402204731   0.9935306494338799   0.1060037257052418   0.42762689203351456   0.46970728033257914   0.48401740617054284   0.08704448053860317   0.23722311528999487   0.4633739612989744   0.16979634100171592   0.503910246185435   0.9528150856841178   0.7167199428912713   0.3776706326398495   0.7274662765794874   0.915223244785385   0.6978702877122946   0.0010962173400467102   0.975126992860913   0.17980736957013616   0.09545491953091863
0.558989525577282   0.9841942804976992   0.8731086148419277   0.4641946793104455   0.5654588761434021   0.8781905547924573   0.4454817228084132   0.9944873989778663   0.08144146997285923   0.7911460742538542   0.20825860751841835   0.531113437678892   0.9116451289711434   0.2872358280684192   0.2554435218343006   0.8143934947876207   0.5339744963312938   0.5597695514889317   0.34022027704891555   0.11652320707532596   0.5328782789912471   0.5846425586280188   0.16041290747877937   0.021068287544407333   0.9738887534139651   0.6004482781303195   0.28730429263685164   0.5568736082339618   0.40842987727056307   0.7222577233378622   0.8418225698284384   0.5623862092560955   0.32698840729770384   0.931111649084008   0.6335639623100201   0.031272771577203526   0.41534327832656054   0.6438758210155888   0.3781204404757195   0.21687927678958288   0.8813687819952668   0.08410626952665706   0.037900163426803996   0.10035606971425692   0.3484905030040197   0.4994637108986383   0.8774872559480246   0.07928778216984958   0.37460174959005454   0.8990154327683187   0.590182963311173   0.5224141739358877   0.9661718723194914   0.1767577094304565   0.7483603934827345   0.9600279646797922   0.6391834650217876   0.2456460603464485   0.1147964311727145   0.9287551931025887   0.22384018669522704   0.6017702393308597   0.736675990696995   0.7118759163130058
0.3424714046999603   0.5176639698042026   0.6987758272701909   0.6115198465987489   0.9939809016959406   0.01820025890556437   0.8212885713221664   0.5322320644288994   0.619379152105886   0.11918482613724568   0.23110560801099336   0.00981789049301161   0.6532072797863946   0.9424271167067891   0.4827452145282588   0.04978992581321934   0.014023814764607009   0.6967810563603407   0.36794878335554426   0.12103473271063059   0.7901836280693799   0.09501081702948094   0.6312727926585493   0.40915881639762475   0.4477122233694197   0.5773468472252783   0.9324969653883584   0.7976389697988757   0.45373132167347907   0.559146588319714   0.111208394066192   0.2654069053699764   0.834352169567593   0.43996176218246824   0.8801027860551986   0.2555890148769648   0.1811448897811984   0.49753464547567905   0.39735757152693985   0.20579908906374547   0.1671210750165914   0.8007535891153384   0.029408788171395566   0.08476435635311487   0.37693744694721143   0.7057427720858575   0.39813599551284623   0.6756055399554901   0.9292252235777918   0.12839592486057916   0.4656390301244879   0.8779665701566144   0.4754939019043127   0.5692493365408652   0.3544306360582959   0.6125596647866379   0.6411417323367197   0.12928757435839697   0.47432785000309724   0.35697064990967314   0.45999684255552126   0.631752928882718   0.0769702784761574   0.1511715608459277
0.29287576753892985   0.8309993397673795   0.04756149030476183   0.06640720449281283   0.9159383205917184   0.12525656768152205   0.6494254947919156   0.3908016645373227   0.9867130970139267   0.9968606428209429   0.1837864646674277   0.5128350943807083   0.511219195109614   0.42761130628007765   0.8293558286091318   0.9002754295940704   0.8700774627728943   0.29832373192168066   0.3550279786060345   0.5433047796843972   0.41008062021737307   0.6665708030389628   0.27805770012987713   0.39213321883846947   0.1172048526784432   0.8355714632715833   0.23049620982511532   0.3257260143456567   0.20126653208672474   0.7103148955900612   0.5810707150331997   0.9349243498083339   0.21455343507279803   0.7134542527691183   0.39728425036577203   0.42208925542762565   0.703334239963184   0.2858429464890407   0.5679284217566403   0.5218138258335553   0.8332567771902897   0.98751921456736   0.21290044315060566   0.9785090461491581   0.4231761569729166   0.32094841152839726   0.9348427430207286   0.5863758273106886   0.3059713042944734   0.485376948256814   0.7043465331956132   0.260649812965032   0.10470477220774864   0.7750620526667528   0.1232758181624135   0.32572546315669804   0.8901513371349506   0.06160779989763441   0.7259915677966414   0.9036362077290724   0.1868170971717666   0.7757648534085937   0.15806314604000124   0.38182238189551704
0.3535603199814769   0.7882456388412337   0.9451627028893955   0.4033133357463589   0.9303841630085603   0.46729722731283646   0.010319959868667045   0.8169375084356703   0.6244128587140869   0.9819202790560225   0.3059734266730538   0.5562876954706383   0.5197080865063383   0.20685822638926976   0.18269760851064035   0.23056223231394024   0.6295567493713877   0.14525042649163533   0.45670604071399884   0.32692602458486786   0.44273965219962114   0.36948557308304164   0.2986428946739976   0.9451036426893509   0.0891793322181442   0.5812399342418079   0.35348019178460205   0.5417903069429919   0.15879516920958386   0.11394270692897142   0.343160231915935   0.7248527985073216   0.5343823104954969   0.1320224278729489   0.03718680524288117   0.16856510303668337   0.014674223989158621   0.9251642014836792   0.8544891967322409   0.9380028707227431   0.3851174746177709   0.7799137749920438   0.397783156018242   0.6110768461378753   0.9423778224181498   0.4104282019090022   0.09914026134424435   0.6659732034485244   0.8531984902000056   0.8291882676671943   0.7456600695596423   0.12418289650553248   0.6944033209904218   0.7152455607382229   0.4024998376437073   0.39933009799821084   0.16002101049492484   0.5832231328652739   0.36531303240082613   0.23076499496152747   0.1453467865057662   0.6580589313815948   0.5108238356685852   0.29276212423878434
0.7602293118879953   0.8781451563895509   0.11304067965034333   0.6816852781009092   0.8178514894698454   0.4677169544805488   0.013900418306098982   0.015712074652384726   0.9646529992698398   0.6385286868133545   0.2682403487464567   0.8915291781468523   0.2702496782794181   0.9232831260751316   0.8657405111027494   0.4921990801486414   0.11022866778449326   0.34005999320985764   0.5004274787019233   0.2614340851871139   0.9648818812787271   0.6820010618282628   0.9896036430333379   0.9686719609483295   0.20465256939073176   0.8038559054387119   0.8765629633829946   0.28698668284742046   0.3868010799208863   0.3361389509581631   0.8626625450768957   0.27127460819503574   0.4221480806510464   0.6976102641448086   0.5944221963304389   0.3797454300481835   0.15189840237162833   0.774327138069677   0.7286816852276896   0.8875463498995421   0.04166973458713506   0.4342671448598194   0.22825420652576633   0.6261122647124282   0.076787853308408   0.7522660830315565   0.2386505634924284   0.6574403037640986   0.8721352839176763   0.9484101775928447   0.3620876001094338   0.37045362091667816   0.48533420399678995   0.6122712266346816   0.4994250550325382   0.09917901272164241   0.0631861233457435   0.914660962489873   0.9050028587020993   0.7194335826734589   0.9112877209741151   0.14033382442019599   0.17632117347440968   0.8318872327739169
0.8696179863869801   0.7060666795603766   0.9480669669486433   0.20577496806148868   0.7928301330785721   0.9538005965288201   0.7094164034562149   0.5483346642973901   0.9206948491608958   0.005390418935975343   0.3473288033467811   0.17788104338071198   0.43536064516410594   0.3931191923012937   0.847903748314243   0.07870203065906956   0.3721745218183624   0.4784582298114207   0.9429008896121437   0.35926844798561064   0.46088680084424727   0.33812440539122474   0.766579716137734   0.5273812152116938   0.5912688144572672   0.6320577258308481   0.8185127491890907   0.3216062471502051   0.7984386813786951   0.6782571293020281   0.10909634573287579   0.7732715828528149   0.8777438322177992   0.6728667103660527   0.7617675423860947   0.5953905394721031   0.4423831870536933   0.279747518064759   0.9138637940718517   0.5166885088130334   0.07020866523533084   0.8012892882533383   0.970962904459708   0.15742006082742283   0.6093218643910836   0.4631648828621136   0.20438318832197397   0.630038845615729   0.01805304993381639   0.8311071570312655   0.38587043913288327   0.30843259846552395   0.21961436855512131   0.1528500277292374   0.27677409340000747   0.5351610156127089   0.34187053633732206   0.47998331736318467   0.5150065510139128   0.9397704761406059   0.8994873492836288   0.20023579929842567   0.6011427569420611   0.4230819673275725
0.829278684048298   0.3989465110450874   0.6301798524823531   0.2656619065001496   0.2199568196572144   0.9357816281829738   0.4257966641603791   0.6356230608844206   0.201903769723398   0.10467447115170833   0.03992622502749585   0.32719046241889665   0.9822894011682767   0.951824443422471   0.7631521316274884   0.7920294468061877   0.6404188648309546   0.4718411260592863   0.24814558061357558   0.8522589706655818   0.7409315155473258   0.27160532676086063   0.6470028236715145   0.42917700333800934   0.9116528314990279   0.8726588157157733   0.01682297118916142   0.16351509683785972   0.6916960118418135   0.9368771875327995   0.5910263070287823   0.5278920359534391   0.48979224211841543   0.8322027163810911   0.5511000820012865   0.20070157353454252   0.5075028409501388   0.8803782729586203   0.7879479503737981   0.4086721267283548   0.8670839761191842   0.40853714689933396   0.5398023697602226   0.556413156062773   0.12615246057185836   0.13693182013847333   0.892799546088708   0.12723615272476366   0.21449962907283052   0.2642730044227001   0.8759765748995466   0.9637210558869039   0.5228036172310171   0.3273958168899006   0.2849502678707643   0.43582901993346473   0.03301137511260161   0.49519310050880944   0.7338501858694778   0.23512744639892225   0.5255085341624628   0.6148148275501892   0.9459022354956798   0.8264553196705675
0.6584245580432787   0.20627768065085528   0.4060998657354572   0.2700421636077945   0.5322720974714203   0.06934586051238195   0.5133003196467492   0.14280601088303083   0.31777246839858975   0.8050728560896819   0.6373237447472027   0.1790849549961269   0.7949688511675727   0.47767703919978133   0.3523734768764384   0.7432559350626622   0.7619574760549711   0.982483938690972   0.6185232910069606   0.5081284886637399   0.23644894189250826   0.3676691111407827   0.6726210555112808   0.6816731689931724   0.5780243838492296   0.1613914304899274   0.2665211897758236   0.411631005385378   0.045752286377809266   0.09204556997754545   0.7532208701290745   0.26882499450234715   0.7279798179792195   0.28697271388786355   0.1158971253818718   0.08974003950622025   0.9330109668116467   0.8092956746880823   0.7635236485054334   0.3464841044435581   0.1710534907566757   0.8268117359971103   0.14500035749847287   0.8383556157798182   0.9346045488641674   0.4591426248563276   0.472379301987192   0.15668244678664578   0.3565801650149379   0.29775119436640024   0.20585811221136838   0.7450514414012678   0.31082787863712863   0.20570562438885476   0.45263724208229394   0.47622644689892063   0.5828480606579092   0.9187329105009912   0.33674011670042214   0.3864864073927004   0.6498370938462623   0.10943723581290897   0.5732164681949887   0.04000230294914229
0.4787836030895866   0.28262549981579865   0.42821611069651583   0.20164668716932407   0.5441790542254191   0.823482874959471   0.9558368087093237   0.04496424038267832   0.18759888921048126   0.5257316805930707   0.7499786964979555   0.29991279898141054   0.8767710105733526   0.32002605620421604   0.29734145441566145   0.8236863520824899   0.2939229499154435   0.40129314570322483   0.9606013377152394   0.4371999446897895   0.6440858560691812   0.29185590989031585   0.38738486952025064   0.3971976417406472   0.16530225297959455   0.009230410074517217   0.9591687588237349   0.19555095457132313   0.6211231987541754   0.18574753511504621   0.003331950114411058   0.1505867141886448   0.43352430954369414   0.6600158545219754   0.25335325361645566   0.8506739152072342   0.5567532989703415   0.3399897983177594   0.9560117992007942   0.026987563124744388   0.262830349054898   0.9386966526145346   0.9954104614855548   0.5897876184349549   0.6187444929857168   0.6468407427242188   0.6080255919653041   0.1925899766943077   0.4534422400061222   0.6376103326497016   0.6488568331415693   0.9970390221229846   0.8323190412519469   0.4518627975346553   0.6455248830271583   0.8464523079343398   0.3987947317082527   0.7918469430126799   0.3921716294107026   0.9957783927271054   0.8420414327379112   0.45185714469492044   0.43615983020990845   0.9687908296023611
0.5792110836830132   0.5131604920803858   0.4407493687243536   0.3790032111674062   0.9604665906972965   0.8663197493561672   0.8327237767590495   0.18641323447309852   0.5070243506911742   0.2287094167064656   0.18386694361748018   0.18937421235011395   0.6747053094392274   0.7768466191718103   0.538342060590322   0.3429219044157742   0.2759105777309747   0.9849996761591304   0.14617043117961934   0.34714351168866875   0.43386914499306345   0.53314253146421   0.7100106009697109   0.3783526820863077   0.8546580613100502   0.019982039383824122   0.26926123224535725   0.9993494709189015   0.8941914706127537   0.153662290027657   0.4365374554863078   0.8129362364458029   0.3871671199215795   0.9249528733211914   0.2526705118688276   0.623562024095689   0.712461810482352   0.14810625414938106   0.7143284512785056   0.28064011967991476   0.43655123275137736   0.1631065779902506   0.5681580200988863   0.933496607991246   0.0026820877583139174   0.6299640465260407   0.8581474191291755   0.5551439259049383   0.14802402644826373   0.6099820071422165   0.5888861868838181   0.5557944549860369   0.25383255583551   0.4563197171145595   0.15234873139751035   0.7428582185402339   0.8666654359139305   0.5313668437933682   0.8996782195286828   0.119296194444545   0.15420362543157848   0.38326058964398707   0.18534976825017707   0.8386560747646302
0.7176523926802011   0.2201540116537365   0.6171917481512907   0.9051594667733842   0.7149703049218872   0.5901899651276958   0.7590443290221154   0.3500155408684459   0.5669462784736234   0.9802079579854794   0.1701581421382972   0.7942210858824089   0.31311372263811343   0.5238882408709199   0.017809410740786836   0.051362867342174996   0.4464482867241829   0.9925213970775517   0.1181311912121041   0.93206667289763   0.29224466129260446   0.6092608074335647   0.932781422961927   0.09341059813299973   0.5745922686124033   0.3891067957798282   0.31558967481063627   0.1882511313596155   0.8596219636905161   0.7989168306521324   0.556545345788521   0.8382355904911696   0.2926756852168927   0.8187088726666529   0.3863872036502238   0.044014504608760635   0.9795619625787793   0.29482063179573303   0.36857779290943693   0.9926516372665857   0.5331136758545963   0.3022992347181813   0.25044660169733285   0.060584964368955656   0.24086901456199192   0.6930384272846166   0.3176651787354058   0.9671743662359559   0.6662767459495886   0.3039316315047884   0.0020755039247695173   0.7789232348763404   0.8066547822590724   0.505014800852656   0.4455301581362486   0.9406876443851708   0.5139790970421797   0.6863059281860031   0.05914295448602479   0.8966731397764102   0.5344171344634004   0.3914852963902701   0.6905651615765879   0.9040215025098246
0.0013034586088040998   0.08918606167208878   0.440118559879255   0.8434365381408689   0.7604344440468122   0.3961476343874722   0.12245338114384921   0.876262171904913   0.0941576980972236   0.09221600288268376   0.1203778772190797   0.09733893702857253   0.2875029158381512   0.5872012020300277   0.6748477190828311   0.15665129264340172   0.7735238187959714   0.9008952738440246   0.6157047645968063   0.2599781528669915   0.239106684332571   0.5094099774537545   0.9251396030202185   0.35595665035716695   0.23780322572376691   0.4202239157816657   0.4850210431409635   0.5125201122162981   0.47736878167695473   0.02407628139419353   0.36256766199711427   0.636257940311385   0.3832110835797311   0.9318602785115098   0.24218978477803457   0.5389190032828125   0.09570816774157995   0.3446590764814821   0.5673420656952034   0.38226771063941084   0.3221843489456085   0.4437638026374575   0.9516373010983971   0.12228955777241933   0.08307766461303746   0.934353825183703   0.02649769807817857   0.7663329074152524   0.8452744388892706   0.5141299094020373   0.5414766549372151   0.2538127951989543   0.36790565721231583   0.4900536280078438   0.17890899294010082   0.6175548548875692   0.9846945736325847   0.558193349496334   0.9367192081620662   0.07863585160475663   0.8889864058910047   0.21353427301485198   0.3693771424668629   0.6963681409653458
0.5668020569453962   0.7697704703773944   0.41773984136846576   0.5740785831929265   0.4837243923323588   0.8354166451936914   0.3912421432902872   0.8077456757776741   0.6384499534430882   0.32128673579165407   0.8497654883530721   0.5539328805787198   0.2705442962307724   0.8312331077838102   0.6708564954129713   0.9363780256911507   0.28584972259818775   0.2730397582874762   0.734137287250905   0.857742174086394   0.396863316707183   0.05950548527262423   0.3647601447840422   0.16137403312104823   0.8300612597617868   0.2897350148952298   0.9470203034155764   0.5872954499281218   0.346336867429428   0.4543183697015384   0.5557781601252891   0.7795497741504477   0.7078869139863397   0.13303163390988432   0.706012671772217   0.22561689357172784   0.4373426177555673   0.30179852612607405   0.035156176359245776   0.28923886788057723   0.15149289515737954   0.028758767838597876   0.3010188891083408   0.4314966937941832   0.7546295784501965   0.9692532825659737   0.9362587443242986   0.27012266067313495   0.9245683186884097   0.6795182676707439   0.9892384409087223   0.6828272107450132   0.5782314512589818   0.22519989796920548   0.43346028078343307   0.9032774365945655   0.870344537272642   0.09216826405932114   0.727447609011216   0.6776605430228376   0.43300191951707473   0.790369737933247   0.6922914326519702   0.38842167514226045
0.2815090243596952   0.7616109700946492   0.39127254354362945   0.9569249813480772   0.5268794459094986   0.7923576875286755   0.45501379921933083   0.6868023206749423   0.6023111272210889   0.1128394198579317   0.4657753583106086   0.0039751099299290965   0.02407967596210711   0.8876395218887262   0.03231507752717556   0.10069767333536359   0.15373513868946506   0.7954712578294051   0.3048674685159595   0.42303713031252593   0.7207332191723903   0.0051015198961580155   0.6125760358639893   0.03461545517026549   0.4392241948126951   0.24349054980150883   0.22130349232035987   0.07769047382218824   0.9123447489031964   0.4511328622728333   0.766289693101029   0.39088815314724595   0.3100336216821075   0.3382934424149016   0.3005143347904204   0.38691304321731684   0.28595394572000044   0.45065392052617537   0.26819925726324484   0.2862153698819533   0.13221880703053535   0.6551826626967703   0.9633317887472853   0.8631782395694273   0.41148558785814504   0.6500811428006122   0.35075575288329597   0.8285627843991619   0.97226139304545   0.40659059299910344   0.1294522605629361   0.7508723105769736   0.05991664414225353   0.9554577307262702   0.36316256746190706   0.35998415742972767   0.749883022460146   0.6171642883113686   0.0626482326714867   0.9730711142124108   0.4639290767401456   0.1665103677851932   0.7944489754082419   0.6868557443304575
0.33171026970961026   0.511327705088423   0.8311171866609566   0.8236775047610302   0.9202246818514652   0.8612465622878106   0.4803614337776606   0.9951147203618683   0.9479632888060152   0.45465596928870716   0.35090917321472453   0.24424240978489467   0.8880466446637617   0.499198238562437   0.9877466057528175   0.884258252355167   0.13816362220361567   0.8820339502510685   0.9250983730813308   0.9111871381427562   0.6742345454634701   0.7155235824658752   0.1306493976730889   0.22433139381229875   0.34252427575385985   0.20419587737745235   0.2995322110121323   0.4006538890512686   0.4222995939023947   0.3429493150896417   0.8191707772344716   0.4055391686894003   0.4743363050963794   0.8882933458009346   0.46826160401974715   0.16129675890450565   0.5862896604326178   0.38909510723849755   0.48051499826692967   0.2770385065493386   0.4481260382290021   0.5070611569874292   0.555416625185599   0.3658513684065824   0.773891492765532   0.7915375745215538   0.42476722751251006   0.14151997459428362   0.4313672170116722   0.5873416971441016   0.12523501650037774   0.740866085543015   0.009067623109277504   0.2443923820544598   0.3060642392659061   0.3353269168536147   0.5347313180128981   0.35609903625352524   0.8378026352461589   0.17403015794910906   0.9484416575802803   0.9670039290150277   0.3572876369792293   0.8969916513997704
0.5003156193512782   0.45994277202759865   0.8018710117936303   0.531140282993188   0.7264241265857462   0.6684051975060448   0.3771037842811203   0.38962030839890444   0.29505690957407404   0.08106350036194324   0.2518687677807425   0.6487542228558895   0.28598928646479654   0.8366711183074834   0.9458045285148364   0.31342730600227475   0.7512579684518985   0.4805720820539582   0.10800189326867748   0.13939714805316566   0.8028163108716182   0.5135681530389304   0.7507142562894482   0.24240549665339522   0.30250069152034   0.05362538101133184   0.9488432444958179   0.7112652136602071   0.5760765649345938   0.3852201835052871   0.5717394602146976   0.3216449052613027   0.2810196553605197   0.3041566831433438   0.3198706924339551   0.6728906824054133   0.9950303688957232   0.4674855648358604   0.3740661639191187   0.3594633764031385   0.2437724004438247   0.9869134827819022   0.2660642706504412   0.22006622834997283   0.44095608957220656   0.4733453297429718   0.5153500143609929   0.9776607316965776   0.13845539805186657   0.4197199487316399   0.5665067698651751   0.26639551803637046   0.5623788331172728   0.03449976522635284   0.9947673096504774   0.9447506127750678   0.2813591777567531   0.730343082083009   0.6748966172165224   0.27185993036965456   0.2863288088610299   0.2628575172471486   0.30083045329740377   0.9123965539665161
0.04255640841720522   0.2759440344652464   0.034766182646962566   0.6923303256165432   0.6016003188449986   0.8025987047222747   0.5194161682859696   0.7146695939199657   0.4631449207931321   0.3828787559906347   0.9529093984207946   0.44827407588359514   0.9007660876758593   0.34837899076428186   0.958142088770317   0.5035234631085274   0.6194069099191062   0.6180359086812729   0.28324547155379465   0.2316635327388728   0.3330781010580762   0.3551783914341243   0.9824150182563909   0.31926697877235677   0.290521692640871   0.07923435696887787   0.9476488356094284   0.6269366531558135   0.6889213737958724   0.27663565224660325   0.42823266732345877   0.9122670592358479   0.22577645300274024   0.8937568962559685   0.4753232689026642   0.46399298335225275   0.325010365326881   0.5453779054916866   0.5171811801323472   0.9604695202437254   0.7056034554077748   0.9273419968104137   0.2339357085785525   0.7288059875048526   0.3725253543496986   0.5721636053762895   0.25152069032216157   0.4095390087324958   0.08200366170882753   0.4929292484074116   0.3038718547127332   0.7826023555766823   0.3930822879129552   0.21629359616080837   0.8756391873892745   0.8703352963408344   0.16730583491021492   0.32253669990483985   0.40031591848661024   0.40634231298858164   0.8422954695833339   0.7771587944131533   0.883134738354263   0.4458727927448562
0.13669201417555915   0.8498167976027395   0.6491990297757106   0.7170668052400035   0.7641666598258606   0.2776531922264501   0.397678339453549   0.3075277965075077   0.6821629981170331   0.7847239438190384   0.09380648474081582   0.5249254409308254   0.2890807102040779   0.5684303476582301   0.21816729735154136   0.6545901445899911   0.12177487529386297   0.24589364775339023   0.8178513788649311   0.24824783160140942   0.27947940571052904   0.46873485334023696   0.934716640510668   0.8023750388565533   0.14278739153496986   0.6189180557374975   0.2855176107349574   0.08530823361654961   0.37862073170910926   0.34126486351104734   0.8878392712814084   0.7777804371090419   0.6964577335920762   0.5565409196920089   0.7940327865405925   0.25285499617821644   0.4073770233879983   0.9881105720337788   0.5758654891890512   0.5982648515882254   0.2856021480941353   0.7422169242803885   0.7580141103241201   0.35001701998681595   0.0061227423836063034   0.27348207094015164   0.8232974698134521   0.5476419811302627   0.8633353508486364   0.6545640152026542   0.5377798590784947   0.46233374751371314   0.4847146191395272   0.3132991516916068   0.6499405877970863   0.6845533104046713   0.788256885547451   0.7567582319995979   0.8559078012564937   0.4316983142264548   0.3808798621594527   0.7686476599658191   0.2800423120674425   0.8334334626382295
0.09527771406531738   0.02643073568543053   0.5220282017433224   0.4834164426514135   0.08915497168171108   0.7529486647452789   0.6987307319298703   0.9357744615211507   0.22581962083307464   0.09838464954262473   0.16095087285137571   0.4734407140074376   0.7411050016935474   0.7850854978510179   0.5110102850542895   0.7888874036027663   0.9528481161460964   0.028327265851419998   0.6551024837977958   0.3571890893763115   0.5719682539866437   0.2596796058856009   0.3750601717303532   0.5237556267380821   0.4766905399213264   0.23324887020017035   0.8530319699870308   0.04033918408666859   0.3875355682396153   0.48030020545489144   0.15430123805716045   0.10456472256551787   0.1617159474065407   0.3819155559122667   0.9933503652057848   0.6311240085580803   0.42061094571299323   0.5968300580612488   0.4823400801514953   0.8422366049553139   0.4677628295668968   0.5685027922098288   0.8272375963536995   0.48504751557900244   0.895794575580253   0.3088231863242279   0.4521774246233463   0.9612918888409203   0.4191040356589266   0.07557431612405756   0.5991454546363155   0.9209527047542517   0.03156846741931128   0.5952741106691661   0.444844216579155   0.8163879821887339   0.8698525200127706   0.2133585547568994   0.4514938513733703   0.18526397363065364   0.44924157429977735   0.6165284966956506   0.969153771221875   0.3430273686753397
0.9814787447328805   0.04802570448582178   0.14191617486817543   0.8579798530963373   0.08568416915262757   0.7392025181615939   0.6897387502448291   0.896687964255417   0.6665801334937009   0.6636282020375363   0.0905932956085136   0.9757352595011651   0.6350116660743896   0.06835409136837017   0.6457490790293585   0.15934727731243123   0.765159146061619   0.8549955366114708   0.1942552276559883   0.9740833036817775   0.31591757176184176   0.2384670399158202   0.2251014564341133   0.6310559350064379   0.33443882702896116   0.19044133542999842   0.0831852815659379   0.7730760819101006   0.2487546578763336   0.45123881726840454   0.3934465313211088   0.8763881176546836   0.5821745243826326   0.7876106152308683   0.3028532357125952   0.9006528581535185   0.947162858308243   0.719256523862498   0.6571041566832366   0.7413055808410873   0.18200371224662387   0.8642609872510273   0.46284892902724833   0.7672222771593097   0.8660861404847822   0.6257939473352071   0.23774747259313503   0.13616634215287182   0.531647313455821   0.4353526119052087   0.15456219102719712   0.36309026024277125   0.28289265557948734   0.9841137946368042   0.7611156597060883   0.4867021425880876   0.7007181311968547   0.1965031794059359   0.45826242399349315   0.586049284434569   0.7535552728886118   0.47724665554343787   0.8011582673102565   0.8447437035934818
0.5715515606419879   0.6129856682924105   0.3383093382830082   0.07752142643417212   0.7054654201572058   0.9871917209572034   0.10056186568987313   0.9413550842813003   0.17381810670138484   0.5518391090519947   0.945999674662676   0.5782648240385291   0.8909254511218975   0.5677253144151906   0.18488401495658768   0.09156268145044141   0.19020731992504275   0.3712221350092547   0.7266215909630945   0.5055133970158723   0.436652047036431   0.8939754794658169   0.925463323652838   0.6607696934223904   0.865100486394443   0.2809898111734063   0.5871539853698299   0.5832482669882184   0.1596350662372373   0.29379809021620285   0.48659211967995675   0.6418931827069181   0.9858169595358525   0.7419589811642081   0.5405924450172808   0.06362835866838908   0.094891508413955   0.17423366674901744   0.3557084300606931   0.9720656772179477   0.9046841884889122   0.8030115317397627   0.6290868390975985   0.46655228020207534   0.46803214145248123   0.9090360522739458   0.7036235154447605   0.8057825867796848   0.6029316550580381   0.6280462411005395   0.11646953007493062   0.22253431979146646   0.44329658882080086   0.3342481508843367   0.6298774103949739   0.5806411370845483   0.4574796292849484   0.5922891697201286   0.08928496537769315   0.5170127784161593   0.3625881208709934   0.41805550297111116   0.7335765353170001   0.5449471011982117
0.45790393238208116   0.6150439712313485   0.10448969621940157   0.0783948209961363   0.9898717909295999   0.7060079189574026   0.4008661807746411   0.2726122342164515   0.38694013587156173   0.07796167785686309   0.2843966506997105   0.050077914424985014   0.9436435470507608   0.7437135269725265   0.6545192403047366   0.46943677734043665   0.48616391776581247   0.15142435725239783   0.5652342749270435   0.9524239989242773   0.12357579689481905   0.7333688542812866   0.8316577396100433   0.4074768977260657   0.6656718645127379   0.11832488304993823   0.7271680433906418   0.32908207672992945   0.675800073583138   0.4123169640925356   0.3263018626160007   0.05646984251347796   0.28885993771157625   0.3343552862356725   0.04190521191629023   0.0063919280884929455   0.3452163906608154   0.5906417592631461   0.38738597161155364   0.5369551507480563   0.859052472895003   0.43921740201074827   0.8221516966845102   0.5845311518237789   0.7354766760001838   0.7058485477294616   0.9904939570744669   0.1770542540977132   0.06980481148744598   0.5875236646795233   0.2633259136838251   0.8479721773677837   0.394004737904308   0.17520670058698776   0.9370240510678244   0.7915023348543058   0.10514480019273172   0.8408514143513153   0.8951188391515341   0.7851104067658129   0.7599284095319163   0.2502096550881691   0.5077328675399805   0.24815525601775656
0.9008759366369133   0.8109922530774208   0.6855811708554703   0.6636241041939777   0.16539926063672947   0.10514370534795923   0.6950872137810035   0.48656985009626447   0.09559444914928347   0.5176200406684358   0.4317613000971784   0.6385976727284807   0.7015897112449755   0.3424133400814481   0.49473724902935406   0.8470953378741749   0.5964449110522437   0.5015619257301329   0.5996184098778199   0.06198493110836203   0.8365165015203275   0.25135227064196375   0.09188554233783942   0.8138296750906054   0.9356405648834141   0.4403600175645429   0.40630437148236914   0.1502055708966278   0.7702413042466847   0.3352163122165837   0.7112171577013656   0.6636357208003634   0.6746468550974012   0.8175962715481478   0.2794558576041873   0.02503804807188268   0.9730571438524257   0.4751829314666997   0.7847186085748332   0.1779427101977078   0.3766122328001819   0.9736210057365668   0.18510019869701333   0.11595777908934576   0.5400957312798544   0.7222687350946031   0.0932146563591739   0.3021281039987403   0.6044551663964404   0.28190871753006014   0.6869102848768048   0.15192253310211248   0.8342138621497557   0.9466924053134764   0.9756931271754391   0.48828681230174914   0.1595670070523545   0.12909613376532864   0.6962372695712519   0.46324876422986644   0.1865098631999288   0.6539132022986289   0.9115186609964185   0.28530605403215864
0.8098976303997468   0.6802921965620621   0.7264184622994052   0.16934827494281288   0.2698018991198924   0.958023461467459   0.6332038059402314   0.8672201709440726   0.665346732723452   0.6761147439373989   0.9462935210634266   0.7152976378419601   0.8311328705736964   0.7294223386239224   0.9706003938879875   0.22701082554021096   0.671565863521342   0.6003262048585938   0.27436312431673565   0.7637620613103445   0.4850560003214131   0.9464130025599649   0.36284446332031706   0.4784560072781859   0.6751583699216662   0.2661208059979028   0.6364260010209117   0.309107732335373   0.40535647080177384   0.3080973445304438   0.003222195080680423   0.4418875613913004   0.7400097380783218   0.631982600593045   0.05692867401725385   0.7265899235493404   0.9088768675046254   0.9025602619691225   0.08632828012926638   0.49957909800912936   0.2373110039832835   0.3022340571105288   0.8119651558125307   0.7358170366987848   0.7522550036618704   0.35582105455056395   0.4491206924922137   0.25736102942059896   0.0770966337402041   0.08970024855266116   0.8126946914713019   0.948253297085226   0.6717401629384302   0.7816029040222173   0.8094724963906215   0.5063657356939255   0.9317304248601085   0.1496203034291724   0.7525438223733677   0.7797758121445852   0.022853557355483035   0.24706004146004984   0.6662155422441013   0.2801967141354558
0.7855425533721996   0.944825984349521   0.8542503864315705   0.5443796774366709   0.03328754971032918   0.5890049297989571   0.4051296939393568   0.287018648016072   0.9561909159701251   0.4993046812462959   0.5924350024680549   0.33876535093084603   0.2844507530316948   0.7177017772240786   0.7829625060774333   0.8323996152369205   0.3527203281715864   0.5680814737949061   0.0304186837040657   0.05262380309233529   0.3298667708161034   0.3210214323348563   0.3642031414599644   0.7724270889568795   0.5443242174439038   0.3761954479853353   0.5099527550283939   0.2280474115202085   0.5110366677335747   0.7871905181863782   0.10482306108903709   0.9410287635041364   0.5548457517634495   0.28788583694008224   0.5123880586209822   0.6022634125732904   0.2703949987317547   0.5701840597160037   0.7294255525435489   0.76986379733637   0.9176746705601684   0.002102585921097533   0.6990068688394832   0.7172399942440346   0.587807899744065   0.6810811535862412   0.33480372737951875   0.9448129052871552   0.043483682300161135   0.304885705600906   0.8248509723511248   0.7167654937669468   0.5324470145665865   0.5176951874145278   0.7200279112620878   0.7757367302628102   0.9776012628031369   0.2298093504744456   0.20763985264110552   0.1734733176895198   0.7072062640713822   0.6596252907584419   0.47821430009755667   0.40360952035314984
0.7895315935112138   0.6575227048373443   0.7792074312580735   0.6863695261091152   0.20172369376714888   0.9764415512511031   0.44440370387855477   0.7415566208219599   0.15824001146698777   0.6715558456501971   0.61955273152743   0.02479112705501327   0.6257929969004012   0.15386065823566933   0.8995248202653422   0.24905439679220304   0.6481917340972644   0.9240513077612238   0.6918849676242367   0.07558107910268323   0.9409854700258822   0.26442601700278184   0.21367066752667999   0.6719715587495334   0.15145387651466832   0.6069033121654375   0.4344632362686065   0.9856020326404182   0.9497301827475194   0.6304617609143344   0.9900595323900517   0.2440454118184582   0.7914901712805317   0.9589059152641373   0.37050680086262183   0.21925428476344494   0.1656971743801304   0.8050452570284679   0.4709819805972797   0.9701998879712419   0.517505440282866   0.8809939492672442   0.779097012973043   0.8946188088685587   0.5765199702569839   0.6165679322644623   0.565426345446363   0.2226472501190253   0.4250660937423156   0.009664620099024787   0.13096310917775653   0.2370452174786071   0.47533591099479616   0.37920285918469043   0.14090357678770477   0.9929998056601489   0.6838457397142644   0.4202969439205532   0.7703967759250829   0.773745520896704   0.5181485653341341   0.6152516868920853   0.29941479532780324   0.8035456329254621
0.0006431250512680274   0.7342577376248413   0.5203177823547602   0.9089268240569034   0.42412315479428414   0.11768980536037893   0.9548914369083972   0.6862795739378781   0.9990570610519686   0.10802518526135414   0.8239283277306406   0.449234356459271   0.5237211500571725   0.7288223260766638   0.6830247509429359   0.4562345507991221   0.8398754103429079   0.3085253821561105   0.912627975017853   0.6824890299024181   0.32172684500877385   0.6932736952640252   0.6132131796900497   0.878943396976956   0.32108371995750584   0.9590159576391839   0.09289539733528956   0.9700165729200526   0.8969605651632216   0.841326152278805   0.1380039604268924   0.28373699898217447   0.8979035041112531   0.7333009670174508   0.31407563269625177   0.8345026425229035   0.3741823540540807   0.004478640940787163   0.6310508817533159   0.3782680917237814   0.5343069437111727   0.6959532587846766   0.7184229067354629   0.6957790618213633   0.21258009870239886   0.0026795635206514996   0.10520972704541318   0.8168356648444073   0.8914963787448931   0.043663605881467546   0.012314329710123615   0.8468190919243547   0.9945358135816713   0.20233745360266253   0.8743103692832312   0.5630820929421801   0.0966323094704182   0.46903648658521163   0.5602347365869794   0.7285794504192767   0.7224499554163375   0.4645578456444245   0.9291838548336635   0.35031135869549535
0.18814301170516476   0.7686045868597479   0.21076094809820062   0.6545322968741321   0.9755629130027659   0.7659250233390963   0.10555122105278744   0.8376966320297248   0.08406653425787287   0.7222614174576287   0.09323689134266383   0.9908775401053702   0.08953072067620155   0.5199239638549662   0.2189265220594326   0.42779544716318996   0.9928984112057834   0.05088747726975461   0.6586917854724532   0.6992159967439132   0.2704484557894458   0.5863296316253301   0.7295079306387896   0.34890463804841787   0.08230544408428107   0.8177250447655823   0.518746982540589   0.6943723411742858   0.10674253108151519   0.051800021426486015   0.41319576148780157   0.856675709144561   0.02267599682364231   0.32953860396885726   0.31995887014513774   0.8657981690391908   0.9331452761474408   0.809614640113891   0.10103234808570512   0.43800272187600087   0.9402468649416574   0.7587271628441364   0.44234056261325194   0.7387867251320877   0.6697984091522116   0.17239753121880624   0.7128326319744623   0.3898820870836697   0.5874929650679305   0.3546724864532239   0.1940856494338733   0.6955097459093839   0.4807504339864153   0.3028724650267379   0.7808898879460717   0.8388340367648229   0.458074437162773   0.9733338610578807   0.460931017800934   0.9730358677256321   0.5249291610153323   0.16371922094398966   0.3598986697152289   0.5350331458496312
0.5846822960736748   0.4049920580998533   0.9175581071019769   0.7962464207175436   0.9148838869214633   0.23259452688104704   0.20472547512751463   0.4063643336338739   0.32739092185353275   0.8779220404278231   0.010639825693641336   0.7108545877244901   0.8466404878671174   0.5750495754010853   0.22974993774756963   0.8720205509596671   0.38856605070434436   0.6017157143432046   0.7688189199466356   0.898984683234035   0.8636368896890121   0.43799649339921487   0.40892025023140677   0.3639515373844038   0.27895459361533725   0.03300443529936159   0.4913621431294299   0.5677051166668602   0.36407070669387404   0.8004099084183145   0.28663666800191523   0.16134078303298627   0.0366797848403413   0.9224878679904914   0.2759968423082739   0.4504861953084962   0.1900392969732239   0.34743829258940623   0.04624690456070429   0.5784656443488291   0.8014732462688795   0.7457225782462017   0.27742798461406865   0.6794809611147941   0.9378363565798674   0.3077260848469868   0.8685077343826618   0.3155294237303903   0.6588817629645302   0.27472164954762524   0.377145591253232   0.7478243070635301   0.29481105627065607   0.4743117411293107   0.09050892325131676   0.5864835240305438   0.2581312714303148   0.5518238731388192   0.8145120809430428   0.13599732872204762   0.0680919744570909   0.20438558054941303   0.7682651763823386   0.5575316843732185
0.26661872818821136   0.45866300230321133   0.49083719176826995   0.8780507232584244   0.328782371608344   0.1509369174562245   0.6223294573856081   0.5625212995280341   0.6699006086438138   0.8762152679085993   0.24518386613237608   0.814696992464504   0.3750895523731578   0.40190352677928864   0.15467494288105932   0.22821346843396018   0.11695828094284297   0.8500796536404693   0.3401628619380164   0.09221613971191255   0.04886630648575206   0.6456940730910564   0.5718976855556779   0.534684455338694   0.7822475782975407   0.18703107078784503   0.08106049378740794   0.6566337320802696   0.4534652066891967   0.03609415333162052   0.45873103640179985   0.09411243255223549   0.7835645980453828   0.15987888542302123   0.2135471702694238   0.27941544008773145   0.40847504567222503   0.7579753586437326   0.05887222738836449   0.05120197165377131   0.2915167647293821   0.9078957050032632   0.718709365450348   0.9589858319418588   0.24265045824363002   0.26220163191220686   0.14681167989467017   0.42430137660316475   0.46040287994608936   0.0751705611243618   0.06575118610726223   0.7676676445228952   0.006937673256892664   0.039076407792741276   0.6070201497054624   0.6735552119706596   0.22337307521150984   0.87919752236972   0.39347297943603854   0.39413977188292815   0.8148980295392848   0.12122216372598746   0.3346007520476741   0.3429378002291568
0.5233812648099028   0.21332645872272424   0.615891386597326   0.38395196828729805   0.2807308065662727   0.9511248268105174   0.46907970670265586   0.9596505916841334   0.8203279266201834   0.8759542656861556   0.40332852059539365   0.19198294716123823   0.8133902533632906   0.8368778578934143   0.7963083708899312   0.5184277351905786   0.5900171781517808   0.9576803355236942   0.4028353914538927   0.12428796330765045   0.7751191486124961   0.8364581717977068   0.06823463940621864   0.7813501630784936   0.2517378838025933   0.6231317130749826   0.4523432528088926   0.39739819479119554   0.9710070772363206   0.6720068862644651   0.9832635461062368   0.4377476031070622   0.1506791506161373   0.7960526205783096   0.5799350255108431   0.24576465594582397   0.3372888972528466   0.9591747626848953   0.7836266546209119   0.7273369207552454   0.7472717191010657   0.0014944271612009972   0.3807912631670191   0.6030489574475949   0.9721525704885697   0.16503625536349417   0.31255662376080046   0.8216987943691013   0.7204146866859764   0.5419045422885116   0.8602133709519079   0.4243005995779058   0.7494076094496558   0.8698976560240465   0.8769498248456712   0.9865529964708436   0.5987284588335184   0.07384503544573683   0.29701479933482805   0.7407883405250196   0.2614395615806719   0.11467027276084156   0.5133881447139163   0.013451419769774237
0.5141678424796061   0.11317584559964057   0.13259688154689708   0.4104024623221793   0.5420152719910364   0.9481395902361464   0.8200402577860966   0.588703667953078   0.82160058530506   0.40623504794763476   0.9598268868341887   0.16440306837517227   0.07219297585540423   0.5363373919235883   0.08287706198851759   0.1778500719043287   0.47346451702188574   0.46249235647785153   0.7858622626536895   0.4370617313793091   0.21202495544121389   0.34782208371700996   0.27247411793977333   0.4236103116095349   0.6978571129616078   0.2346462381173694   0.13987723639287625   0.013207849287355541   0.15584184097057138   0.28650664788122304   0.3198369786067796   0.42450418133427753   0.3342412556655114   0.8802715999335883   0.3600100917725909   0.26010111295910526   0.2620482798101072   0.34393420800999985   0.27713302978407334   0.08225104105477654   0.7885837627882214   0.8814418515321484   0.4912707671303838   0.6451893096754674   0.5765588073470076   0.5336197678151383   0.21879664919061045   0.22157899806593256   0.8787016943853998   0.29897352969776897   0.07891941279773419   0.20837114877857704   0.7228598534148284   0.01246688181654592   0.7590824341909546   0.7838669674442995   0.388618597749317   0.13219528188295768   0.39907234241836365   0.5237658544851943   0.1265703179392098   0.7882610738729579   0.1219393126342903   0.4415148134304177
0.33798655515098835   0.9068192223408095   0.6306685455039065   0.7963255037549503   0.7614277478039808   0.3731994545256711   0.41187189631329607   0.5747465056890178   0.882726053418581   0.07422592482790218   0.33295248351556184   0.3663753569104407   0.15986620000375262   0.06175904301135626   0.5738700493246073   0.5825083894661411   0.7712476022544357   0.9295637611283986   0.1747977069062437   0.05874253498094689   0.6446772843152259   0.14130268725544076   0.052858394271953386   0.6172277215505292   0.3066907291642375   0.2344834649146313   0.4221898487680469   0.8209022177955788   0.5452629813602566   0.8612840103889602   0.01031795245475082   0.24615571210656115   0.6625369279416756   0.7870580855610579   0.6773654689391889   0.8797803551961204   0.5026707279379231   0.7252990425497017   0.10349541961458164   0.29727196572997927   0.7314231256834874   0.7957352814213031   0.928697712708338   0.2385294307490324   0.08674584136826158   0.6544325941658624   0.8758393184363845   0.6213017091985032   0.7800551122040241   0.41994912925123107   0.4536494696683377   0.8003994914029244   0.2347921308437674   0.5586651188622709   0.4433315172135869   0.5542437792963633   0.5722552029020918   0.7716070333012129   0.765966048274398   0.6744634241002427   0.06958447496416868   0.04630799075151121   0.6624706286598163   0.37719145837026347
0.33816134928068126   0.2505727093302081   0.7337729159514783   0.13866202762123106   0.2514155079124197   0.5961401151643457   0.8579335975150938   0.5173603184227278   0.47136039570839555   0.1761909859131146   0.40428412784675605   0.7169608270198035   0.23656826486462815   0.6175258670508437   0.9609526106331692   0.1627170477234402   0.6643130619625364   0.8459188337496307   0.19498656235877126   0.4882536236231974   0.5947285869983677   0.7996108429981196   0.532515933698955   0.11106216525293394   0.25656723771768647   0.5490381336679114   0.7987430177474767   0.9724001376317029   0.005151729805266782   0.9528980185035658   0.9408094202323829   0.45503981920897507   0.5337913340968712   0.7767070325904512   0.5365252923856269   0.7380789921891716   0.29722306923224306   0.1591811655396075   0.5755726817524577   0.5753619444657314   0.6329100072697066   0.31326233178997676   0.3805861193936864   0.08710832084253398   0.0381814202713389   0.5136514887918572   0.8480701856947315   0.9760461555896001   0.7816141825536524   0.9646133551239457   0.049327167947254745   0.003646017957897154   0.7764624527483857   0.011715336620379952   0.1085177477148718   0.5486061987489221   0.24267111865151444   0.23500830402992876   0.5719924553292449   0.8105272065597505   0.9454480494192714   0.07582713849032127   0.9964197735767872   0.23516526209401908
0.31253804214956477   0.7625648067003445   0.6158336541831008   0.1480569412514851   0.27435662187822585   0.2489133179084873   0.7677634684883693   0.17201078566188507   0.49274243932457346   0.28429996278454156   0.7184363005411145   0.16836476770398792   0.7162799865761877   0.2725846261641616   0.6099185528262427   0.6197585689550659   0.4736088679246733   0.037576322134232835   0.037926097496997865   0.8092313623953153   0.5281608185054019   0.9617491836439116   0.041506323920210676   0.5740661003012962   0.21562277635583713   0.19918437694356705   0.42567266973710993   0.4260091590498111   0.9412661544776113   0.9502710590350798   0.6579092012487406   0.253998373387926   0.44852371515303785   0.6659710962505382   0.939472900707626   0.08563360568393812   0.73224372857685   0.3933864700863766   0.32955434788138327   0.46587503672887226   0.2586348606521767   0.3558101479521438   0.2916282503843854   0.656643674333557   0.7304740421467748   0.3940609643082322   0.25012192646417475   0.08257757403226071   0.5148512657909377   0.19487658736466512   0.8244492567270648   0.6565684149824496   0.5735851113133265   0.24460552832958538   0.1665400554783242   0.40257004159452353   0.12506139616028858   0.5786344320790472   0.22706715477069814   0.3169364359105854   0.39281766758343856   0.18524796199267057   0.8975128068893149   0.8510613991817131
0.1341828069312618   0.8294378140405269   0.6058845565049295   0.19441772484815617   0.403708764784487   0.4353768497322946   0.3557626300407547   0.11184015081589546   0.8888574989935493   0.2405002623676295   0.5313133733136899   0.4552717358334459   0.3152723876802229   0.9958947340380441   0.3647733178353657   0.05270169423892234   0.1902109915199343   0.41726030195899694   0.13770616306466757   0.735765258328337   0.7973933239364958   0.2320123399663264   0.2401933561753527   0.8847038591466238   0.6632105170052339   0.40257452592579956   0.6343087996704232   0.6902861342984676   0.259501752220747   0.9671976761935049   0.27854616962966855   0.5784459834825721   0.3706442532271977   0.7266974138258755   0.7472327963159786   0.12317424764912624   0.05537186554697477   0.7308026797878313   0.3824594784806129   0.0704725534102039   0.8651608740270404   0.3135423778288344   0.24475331541594536   0.334707295081867   0.06776755009054466   0.081530037862508   0.0045599592405926636   0.4500034359352432   0.4045570330853107   0.6789555119367084   0.3702511595701694   0.7597173016367756   0.1450552808645637   0.7117578357432034   0.09170498994050089   0.1812713181542035   0.774411027637366   0.985060421917328   0.34447219362452225   0.058097070505077265   0.7190391620903913   0.2542577421294966   0.9620127151439094   0.9876245170948733
0.8538782880633509   0.9407153643006623   0.717259399727964   0.6529172220130064   0.7861107379728062   0.8591853264381543   0.7126994404873713   0.20291378607776317   0.38155370488749546   0.18022981450144582   0.3424482809172019   0.4431964844409875   0.23649842402293175   0.46847197875824237   0.250743290976701   0.26192516628678403   0.46208739638556573   0.4834115568409144   0.9062710973521787   0.20382809578170677   0.7430482342951744   0.2291538147114178   0.9442583822082694   0.2162035786868334   0.8891699462318237   0.2884384504107556   0.2269989824803054   0.563286356673827   0.10305920825901749   0.42925312397260135   0.514299541992934   0.36037257059606387   0.7215055033715221   0.24902330947115556   0.17185126107573218   0.9171760861550763   0.4850070793485903   0.7805513307129132   0.9211079700990311   0.6552509198682923   0.02291968296302459   0.29713977387199875   0.014836872746852406   0.4514228240865855   0.27987144866785013   0.06798595916058096   0.070578490538583   0.23521924539975214   0.3907015024360265   0.7795475087498254   0.8435795080582776   0.6719328887259252   0.28764229417700904   0.350294384777224   0.32927996606534354   0.3115603181298613   0.566136790805487   0.10127107530606845   0.15742870498961137   0.39438423197478495   0.0811297114568967   0.3207197445931553   0.2363207348905802   0.7391333121064927
0.0582100284938721   0.023579970721156498   0.2214838621437278   0.2877104880199071   0.778338579826022   0.9555940115605756   0.15090537160514478   0.05249124262015496   0.3876370773899954   0.17604650281075016   0.3073258635468672   0.3805583538942298   0.09999478321298641   0.8257521180335261   0.9780458974815237   0.06899803576436855   0.5338579924074994   0.7244810427274577   0.8206171924919123   0.6746138037895836   0.45272828095060275   0.40376129813430245   0.5842964576013321   0.935480491683091   0.3945182524567306   0.3801813274131459   0.3628125954576043   0.6477700036631838   0.6161796726307087   0.4245873158525704   0.2119072238524595   0.5952787610430289   0.22854259524071324   0.24854081304182024   0.9045813603055923   0.21472040714879906   0.12854781202772683   0.4227886950082941   0.9265354628240686   0.1457223713844305   0.5946898196202274   0.6983076522808364   0.10591827033215635   0.47110856759484687   0.1419615386696247   0.29454635414653396   0.5216218127308243   0.535628075911756   0.747443286212894   0.914365026733388   0.15880921727321998   0.887858072248572   0.13126361358218538   0.4897777108808177   0.9469019934207604   0.2925793112055432   0.9027210183414721   0.2412368978389974   0.04232063311516816   0.07785890405674419   0.7741732063137453   0.8184482028307033   0.11578517029109951   0.9321365326723137
0.17948338669351793   0.12014055054986691   0.00986689995894316   0.4610279650774668   0.03752184802389325   0.825594196403333   0.4882450872281189   0.9253998891657108   0.29007856181099917   0.9112291696699448   0.32943586995489893   0.03754181691713875   0.1588149482288138   0.4214514587891272   0.38253387653413845   0.7449625057115955   0.25609392988734164   0.1802145609501298   0.3402132434189703   0.6671036016548514   0.4819207235735963   0.3617663581194265   0.22442807312787078   0.7349670689825376   0.30243733688007834   0.24162580756955956   0.21456117316892762   0.27393910390507087   0.2649154888561851   0.41603161116622667   0.7263160859408088   0.34853921473936   0.9748369270451859   0.5048024414962817   0.3968802159859098   0.31099739782222124   0.8160219788163721   0.08335098270715456   0.014346339451771344   0.5660348921106257   0.5599280489290305   0.9031364217570248   0.674133096032801   0.8989312904557744   0.07800732535543417   0.5413700636375983   0.4497050229049303   0.16396422147323672   0.7755699884753559   0.29974425606803873   0.2351438497360027   0.8900251175681658   0.5106544996191708   0.8837126449018121   0.508827763795194   0.5414859028288058   0.5358175725739848   0.37891020340553033   0.11194754780928418   0.23048850500658458   0.7197955937576127   0.29555922069837576   0.09760120835751283   0.6644536128959588
0.15986754482858223   0.39242279894135096   0.42346811232471177   0.7655223224401845   0.08186021947314805   0.8510527353037527   0.9737630894197815   0.6015581009669477   0.30629023099779223   0.5513084792357139   0.7386192396837788   0.7115329833987819   0.7956357313786215   0.6675958343339019   0.22979147588858484   0.170047080569976   0.2598181588046367   0.2886856309283715   0.11784392807930065   0.9395585755633914   0.5400225650470241   0.9931264102299958   0.020242719721787813   0.27510496266743256   0.3801550202184418   0.6007036112886448   0.596774607397076   0.5095826402272481   0.29829480074529374   0.7496508759848921   0.6230115179772946   0.9080245392603004   0.9920045697475015   0.19834239674917817   0.8843922782935157   0.19649155586151854   0.19636883836888   0.5307465624152763   0.6546008024049309   0.02644447529154253   0.9365506795642433   0.24206093148690475   0.5367568743256302   0.08688589972815111   0.39652811451721925   0.24893452125690896   0.5165141546038424   0.8117809370607185   0.016373094298777452   0.6482309099682642   0.9197395472067664   0.30219829683347044   0.7180782935534837   0.898580033983372   0.2967280292294719   0.39417375757317   0.7260737238059822   0.7002376372341939   0.4123357509359561   0.1976822017116515   0.5297048854371023   0.1694910748189176   0.7577349485310252   0.17123772642010898
0.5931542058728589   0.9274301433320129   0.2209780742053949   0.08435182669195786   0.1966260913556397   0.6784956220751039   0.7044639196015524   0.2725708896312393   0.18025299705686224   0.030264712106839738   0.784724372394786   0.9703725927977689   0.4621747035033785   0.1316846781234677   0.4879963431653141   0.5761988352245988   0.7361009796973963   0.4314470408892738   0.07566059222935798   0.37851663351294734   0.20639609426029412   0.2619559660703562   0.3179256436983328   0.20727890709283836   0.6132418883874352   0.33452582273834336   0.09694756949293791   0.1229270804008805   0.4166157970317955   0.6560302006632395   0.3924836498913855   0.8503561907696412   0.23636279997493326   0.6257654885563997   0.6077592774965995   0.8799835979718723   0.7741880964715547   0.494080810432932   0.11976293433128542   0.3037847627472735   0.03808711677415839   0.06263376954365822   0.044102342101927434   0.9252681292343261   0.8316910225138643   0.800677803473302   0.7261766984035947   0.7179892221414877   0.21844913412642908   0.46615198073495867   0.6292291289106567   0.5950621417406072   0.8018333370946336   0.8101217800717192   0.23674547901927123   0.744705950970966   0.5654705371197003   0.18435629151531946   0.6289862015226717   0.8647223529990937   0.7912824406481456   0.6902754810823875   0.5092232671913863   0.5609375902518203
0.7531953238739872   0.6276417115387292   0.46512092508945885   0.6356694610174941   0.921504301360123   0.8269639080654272   0.7389442266858642   0.9176802388760064   0.7030551672336939   0.3608119273304686   0.1097150977752075   0.3226180971353991   0.9012218301390603   0.5506901472587493   0.8729696187559363   0.577912146164433   0.33575129301935996   0.3663338557434299   0.24398341723326455   0.7131897931653393   0.5444688523712143   0.6760583746610425   0.7347601500418782   0.15225220291351896   0.7912735284972272   0.04841666312231326   0.2696392249524194   0.5165827418960248   0.8697692271371043   0.22145275505688605   0.5306949982665552   0.5989025030200185   0.16671405990341037   0.8606408277264175   0.42097990049134765   0.2762844058846194   0.26549222976435005   0.3099506804676681   0.5480102817354113   0.6983722597201865   0.9297409367449901   0.9436168247242382   0.30402686450214683   0.9851824665548472   0.3852720843737757   0.26755845006319573   0.5692667144602686   0.8329302636413283   0.5939985558765485   0.2191417869408825   0.2996274895078492   0.3163475217453034   0.7242293287394442   0.9976890318839965   0.768932491241294   0.717445018725285   0.5575152688360339   0.13704820415757893   0.34795259074994644   0.44116061284066554   0.2920230390716838   0.8270975236899109   0.799942309014535   0.7427883531204791
0.3622821023266937   0.8834806989656726   0.4959154445123882   0.7576058865656319   0.977010017952918   0.6159222489024768   0.9266487300521197   0.9246756229243037   0.3830114620763695   0.39678046196159433   0.6270212405442704   0.6083281011790003   0.6587821333369253   0.3990914300775979   0.8580887493029764   0.8908830824537153   0.10126686450089131   0.262043225920019   0.51013615855303   0.4497224696130498   0.8092438254292075   0.43494570223010814   0.710193849538495   0.7069341164925707   0.44696172310251375   0.5514650032644356   0.2142784050261067   0.9493282299269388   0.4699517051495957   0.9355427543619588   0.28762967497398706   0.024652607002635066   0.08694024307322624   0.5387622924003644   0.6606084344297166   0.4163245058236348   0.42815810973630103   0.1396708623227665   0.8025196851267402   0.5254414233699195   0.3268912452354097   0.8776276364027475   0.2923835265737102   0.07571895375686967   0.5176474198062022   0.44268193417263935   0.5821896770352153   0.368784837264299   0.07068569670368847   0.8912169309082038   0.36791127200910856   0.41945660733736023   0.6007339915540927   0.9556741765462451   0.08028159703512153   0.3948040003347252   0.5137937484808665   0.41691188414588065   0.41967316260540494   0.9784794945110904   0.08563563874456545   0.27724102182311416   0.6171534774786648   0.4530380711411709
0.7587443935091558   0.3996133854203666   0.32476995090495453   0.37731911738430124   0.24109697370295352   0.9569314512477273   0.7425802738697392   0.008534280120002253   0.17041127699926503   0.06571452033952348   0.3746690018606307   0.589077672782642   0.5696772854451723   0.11004034379327844   0.2943874048255092   0.19427367244791685   0.05588353696430583   0.6931284596473978   0.8747142422201042   0.21579417793682648   0.9702478982197403   0.41588743782428367   0.25756076474143946   0.7627561067956555   0.21150350471058463   0.01627405240391701   0.932790813836485   0.3854369894113543   0.9704065310076311   0.05934260115618974   0.1902105399667457   0.37690270929135206   0.7999952540083661   0.9936280808166662   0.815541538106115   0.78782503650871   0.23031796856319378   0.8835877370233878   0.5211541332806059   0.5935513640607932   0.17443443159888797   0.19045927737599003   0.6464398910605016   0.37775718612396675   0.20418653337914758   0.7745718395517064   0.38887912631906213   0.6150010793283112   0.992683028668563   0.7582977871477894   0.4560883124825772   0.22956408991695684   0.0222764976609318   0.6989551859915997   0.2658777725158315   0.8526613806256048   0.2222812436525657   0.7053271051749334   0.4503362344097165   0.06483634411689473   0.9919632750893719   0.8217393681515456   0.9291821011291106   0.47128498005610153
0.8175288434904839   0.6312800907755556   0.282742210068609   0.0935277939321348   0.6133423101113364   0.8567082512238492   0.8938630837495469   0.4785267146038236   0.6206592814427735   0.09841046407605977   0.43777477126696973   0.24896262468686678   0.5983827837818416   0.39945527808446013   0.17189699875113823   0.396301244061262   0.37610154012927594   0.6941281729095268   0.7215607643414218   0.3314648999443673   0.384138265039904   0.8723888047579812   0.7923786632123111   0.8601799198882657   0.5666094215494201   0.2411087139824257   0.5096364531437021   0.766652125956131   0.9532671114380836   0.3844004627585766   0.6157733693941553   0.2881254113523073   0.3326078299953102   0.2859899986825168   0.17799859812718552   0.03916278666544052   0.7342250462134686   0.8865347205980566   0.006101599376047304   0.6428615426041785   0.35812350608419263   0.19240654768852986   0.28454083503462557   0.31139664265981126   0.9739852410442886   0.32001774293054863   0.4921621718223144   0.45121672277154556   0.40737581949486856   0.07890902894812292   0.9825257186786123   0.6845645968154146   0.4541087080567849   0.6945085661895464   0.36675234928445705   0.3964391854631073   0.12150087806147468   0.4085185675070296   0.18875375115727153   0.35727639879766676   0.3872758318480061   0.5219838469089729   0.18265215178122424   0.7144148561934882
0.029152325763813478   0.3295772992204431   0.8981113167465987   0.403018213533677   0.05516708471952487   0.009559556289894444   0.40594914492428424   0.9518014907621315   0.6477912652246564   0.9306505273417716   0.423423426245672   0.26723689394671685   0.19368255716787142   0.23614196115222516   0.05667107696121489   0.8707977084836095   0.07218167910639672   0.8276233936451955   0.8679173258039433   0.5135213096859428   0.6849058472583907   0.3056395467362227   0.6852651740227191   0.7991064534924545   0.6557535214945771   0.9760622475157796   0.7871538572761204   0.3960882399587775   0.6005864367750523   0.9665026912258852   0.3812047123518362   0.444286749196646   0.952795171550396   0.03585216388411362   0.9577812861061642   0.1770498552499292   0.7591126143825245   0.7997102027318884   0.9011102091449493   0.3062521467663197   0.6869309352761278   0.9720868090866929   0.03319288334100598   0.792730837080377   0.002025088017737215   0.6664472623504702   0.34792770931828687   0.9936243835879224   0.3462715665231601   0.6903850148346906   0.5607738520421663   0.5975361436291449   0.7456851297481079   0.7238823236088054   0.1795691396903302   0.15324939443249888   0.7928899581977118   0.6880301597246918   0.22178785358416597   0.9761995391825697   0.03377734381518727   0.8883199569928034   0.32067764443921665   0.66994739241625
0.34684640853905946   0.9162331479061105   0.28748476109821064   0.8772165553358732   0.34482132052132225   0.24978588555564032   0.9395570517799238   0.8835921717479507   0.9985497539981621   0.5594008707209497   0.3787831997377574   0.2860560281188058   0.25286462425005435   0.8355185471121442   0.1992140600474272   0.13280663368630694   0.4599746660523425   0.14748838738745237   0.9774262064632613   0.15660709450373722   0.42619732223715523   0.259168430394649   0.6567485620240446   0.4866597020874872   0.0793509136980958   0.34293528248853844   0.36926380092583394   0.609443146751614   0.7345295931767736   0.09314939693289812   0.4297067491459101   0.7258509750036634   0.7359798391786114   0.5337485262119485   0.050923549408152705   0.4397949468848575   0.4831152149285571   0.6982299790998042   0.8517094893607255   0.3069883131985506   0.023140548876214563   0.5507415917123518   0.8742832828974643   0.15038121869481333   0.5969432266390593   0.29157316131770283   0.21753472087341966   0.6637215166073261   0.5175923129409635   0.9486378788291644   0.8482709199475857   0.05427836985571211   0.78306271976419   0.8554884818962664   0.41856417080167563   0.3284273948520488   0.04708288058557854   0.3217399556843179   0.3676406213935229   0.8886324479671913   0.5639676656570215   0.6235099765845137   0.5159311320327974   0.5816441347686407
0.5408271167808069   0.07276838487216189   0.6416478491353331   0.4312629160738274   0.9438838901417476   0.781195223554459   0.4241131282619135   0.7675413994665012   0.42629157720078403   0.8325573447252946   0.5758422083143278   0.7132630296107891   0.6432288574365941   0.9770688628290283   0.15727803751265215   0.38483563475874033   0.5961459768510156   0.6553289071447104   0.7896374161191292   0.496203186791549   0.032178311193994086   0.03181893056019666   0.2737062840863318   0.9145590520229083   0.4913511944131872   0.9590505456880347   0.6320584349509987   0.4832961359490809   0.5474673042714396   0.17785532213357574   0.20794530668908517   0.7157547364825796   0.12117572707065555   0.3452979774082811   0.6321030983747574   0.002491706871790511   0.47794686963406147   0.36822911457925284   0.4748250608621053   0.6176560721130502   0.8818008927830459   0.7129002074345425   0.685187644742976   0.12145288532150117   0.8496225815890518   0.6810812768743458   0.4114813606566442   0.2068938332985929   0.35827138717586465   0.722030731186311   0.7794229257056455   0.7235976973495121   0.8108040829044251   0.5441754090527353   0.5714776190165604   0.007842960866932381   0.6896283558337695   0.19887743164445418   0.9393745206418029   0.005351253995141869   0.21168148619970803   0.8306483170652014   0.4645494597796977   0.3876951818820917
0.32988059341666215   0.11774810963065885   0.7793618150367216   0.2662422965605905   0.48025801182761035   0.436666832756313   0.36788045438007744   0.0593484632619976   0.12198662465174569   0.714636101570002   0.5884575286744319   0.3357507659124856   0.31118254174732063   0.17046069251726667   0.01697990965787151   0.3279078050455532   0.6215541859135512   0.9715832608728125   0.07760538901606856   0.3225565510504113   0.4098726997138431   0.1409349438076112   0.6130559292363709   0.9348613691683196   0.07999210629718097   0.02318683417695236   0.8336941141996492   0.6686190726077291   0.5997340944695706   0.5865200014206393   0.4658136598195718   0.6092706093457315   0.47774746981782495   0.8718838998506373   0.8773561311451399   0.273519843433246   0.1665649280705043   0.7014232073333707   0.8603762214872684   0.9456120383876928   0.5450107421569531   0.7298399464605582   0.7827708324711998   0.6230554873372814   0.13513804244311003   0.588905002652947   0.169714903234829   0.6881941181689618   0.05514593614592907   0.5657181684759945   0.33602078903517973   0.01957504556123262   0.4554118416763584   0.9791981670553552   0.8702071292156079   0.41030443621550106   0.9776643718585335   0.10731426720471791   0.992850998070468   0.1367845927822551   0.8110994437880291   0.40589105987134727   0.13247477658319956   0.19117255439456235
0.266088701631076   0.6760511134107892   0.34970394411199973   0.5681170670572809   0.13095065918796597   0.08714611075784216   0.17998904087717071   0.8799229488883191   0.0758047230420369   0.5214279422818475   0.843968251841991   0.8603479033270865   0.6203928813656785   0.5422297752264923   0.973761122626383   0.45004346711158544   0.642728509507145   0.4349155080217744   0.9809101245559151   0.31325887432933036   0.8316290657191159   0.029024448150427144   0.8484353479727155   0.122086319934768   0.5655403640880399   0.35297333473963804   0.4987314038607158   0.5539692528774871   0.43458970490007387   0.26582722398179587   0.3187423629835451   0.674046303989168   0.358784981858037   0.7443992816999483   0.4747741111415541   0.8136984006620814   0.7383921004923585   0.20216950647345597   0.5010129885151711   0.36365493355049594   0.09566359098521346   0.7672539984516816   0.520102863959256   0.05039605922116559   0.2640345252660976   0.7382295503012545   0.6716675159865405   0.9283097392863976   0.6984941611780577   0.3852562155616164   0.17293611212582471   0.3743404864089105   0.26390445627798387   0.11942899157982052   0.8541937491422796   0.7002941824197426   0.9051194744199469   0.3750297098798722   0.3794196380007256   0.8865957817576612   0.1667273739275884   0.17286020340641625   0.8784066494855546   0.5229408482071652
0.07106378294237496   0.4056062049547347   0.3583037855262986   0.4725447889859996   0.8070292576762774   0.6673766546534803   0.6866362695397581   0.544235049699602   0.10853509649821964   0.28212043909186385   0.5137001574139334   0.16989456329069152   0.8446306402202358   0.16269144751204334   0.6595064082716537   0.46960038087094896   0.9395111658002889   0.7876617376321711   0.2800867702709282   0.5830045991132877   0.7727837918727005   0.6148015342257548   0.40168012078537363   0.06006375090612255   0.7017200089303255   0.20919532927102014   0.04337633525907505   0.5875189619201229   0.8946907512540482   0.5418186746175399   0.35674006571931693   0.04328391222052087   0.7861556547558285   0.259698235525676   0.8430399083053836   0.8733893489298293   0.9415250145355927   0.09700678801363269   0.18353350003372979   0.40378896805888037   0.0020138487353038334   0.3093450503814616   0.9034467297628016   0.8207843689455926   0.22923005686260337   0.6945435161557068   0.501766608977428   0.7607206180394701   0.5275100479322778   0.4853481868846866   0.45839027371835295   0.17320165611934715   0.6328192966782297   0.9435295122671468   0.10165020799903599   0.12991774389882627   0.8466636419224012   0.6838312767414707   0.25861029969365246   0.25652839496899693   0.9051386273868085   0.586824488727838   0.07507679965992266   0.8527394269101165
0.9031247786515046   0.27747943834637645   0.17163006989712107   0.031955057964523914   0.6738947217889013   0.5829359221906697   0.6698634609196931   0.27123443992505386   0.14638467385662346   0.09758773530598305   0.21147318720134017   0.09803278380570671   0.5135653771783937   0.15405822303883632   0.10982297920230419   0.9681150399068804   0.6669017352559925   0.4702269462973656   0.8512126795086518   0.7115866449378835   0.761763107869184   0.8834024575695276   0.7761358798487291   0.858847218027767   0.8586383292176794   0.6059230192231512   0.6045058099516081   0.8268921600632431   0.18474360742877802   0.022987097032481474   0.9346423490319149   0.5556577201381893   0.03835893357215455   0.9253993617264984   0.7231691618305748   0.4576249363324825   0.5247935563937608   0.7713411386876621   0.6133461826282706   0.48950989642560205   0.8578918211377683   0.30111419239029646   0.7621335031196188   0.7779232514877186   0.09612871326858433   0.4177117348207689   0.9859976232708897   0.9190760334599516   0.237490384050905   0.8117887155976178   0.38149181331928167   0.09218387339670849   0.052746776622127   0.7888016185651363   0.44684946428736677   0.5365261532585193   0.014387843049972447   0.8634022568386378   0.723680302456792   0.07890121692603674   0.48959428665621163   0.09206111815097577   0.11033411982852143   0.5893913205004346
0.6317024655184433   0.7909469257606793   0.3482006167089026   0.8114680690127162   0.535573752249859   0.3732351909399104   0.3622029934380129   0.8923920355527646   0.298083368198954   0.5614464753422926   0.9807111801187312   0.8002081621560561   0.24533659157682697   0.7726448567771563   0.5338617158313644   0.26368200889753685   0.23094874852685454   0.9092425999385185   0.8101814133745724   0.18478079197150007   0.7413544618706429   0.8171814817875428   0.699847293546051   0.5953894714710654   0.1096519963521996   0.026234556026863472   0.3516466768371484   0.7839214024583493   0.5740782441023407   0.6529993650869531   0.9894436833991355   0.8915293669055847   0.2759948759033866   0.09155288974466043   0.00873250328040432   0.0913212047495286   0.030658284326559655   0.31890803296750403   0.4748707874490399   0.8276391958519917   0.7997095357997052   0.4096654330289855   0.6646893740744675   0.6428584038804916   0.05835507392906221   0.5924839512414427   0.9648420805284165   0.04746893240942627   0.9487030775768626   0.5662493952145793   0.613195403691268   0.263547529951077   0.37462483347452197   0.9132500301276262   0.6237517202921325   0.3720181630454923   0.09862995757113535   0.8216971403829658   0.6150192170117282   0.2806969582959637   0.0679716732445757   0.5027891074154618   0.14014842956268836   0.45305776244397195
0.2682621374448706   0.09312367438647622   0.47545905548822087   0.8101993585634802   0.20990706351580837   0.5006397231450335   0.5106169749598044   0.762730426154054   0.2612039859389458   0.9343903279304542   0.8974215712685364   0.499182896202977   0.8865791524644238   0.021140297802827966   0.2736698509764038   0.1271647331574847   0.7879491948932884   0.19944315741986218   0.6586506339646756   0.846467774861521   0.7199775216487128   0.6966540500044004   0.5185022044019872   0.393410012417549   0.4517153842038421   0.6035303756179242   0.043043148913766316   0.5832106538540688   0.24180832068803376   0.10289065247289077   0.5324261739539619   0.8204802277000148   0.980604334749088   0.1685003245424366   0.6350046026854256   0.3212973314970378   0.09402518228466421   0.14736002673960863   0.36133475170902174   0.1941325983395531   0.3060759873913758   0.9479168693197465   0.7026841177443462   0.3476648234780321   0.5860984657426631   0.251262819315346   0.184181913342359   0.954254811060483   0.13438308153882095   0.6477324436974218   0.1411387644285927   0.37104415720641426   0.8925747608507872   0.544841791224531   0.6087125904746308   0.5505639295063995   0.9119704261016992   0.3763414666820944   0.9737079877892052   0.2292665980093617   0.817945243817035   0.22898143994248576   0.6123732360801835   0.03513399966980859
0.5118692564256592   0.2810645706227393   0.9096891183358373   0.6874691761917765   0.9257707906829962   0.029801751307393314   0.7255072049934783   0.7332143651312935   0.7913877091441752   0.38206930760997154   0.5843684405648856   0.36217020792487914   0.898812948293388   0.8372275163854406   0.9756558500902548   0.8116062784184797   0.9868425221916888   0.4608860497033461   0.0019478623010495666   0.582339680409118   0.1688972783746538   0.2319046097608604   0.3895746262208661   0.5472056807393093   0.6570280219489946   0.9508400391381211   0.4798855078850288   0.8597365045475329   0.7312572312659984   0.9210382878307277   0.7543783028915505   0.12652213941623947   0.9398695221218233   0.5389689802207562   0.17000986232666493   0.7643519314913604   0.04105657382843528   0.7017414638353157   0.1943540122364101   0.9527456530728807   0.05421405163674649   0.2408554141319695   0.19240614993536057   0.37040597266376274   0.8853167732620927   0.008950804371109131   0.8028315237144945   0.8232002919244534   0.22828875131309811   0.05811076523298807   0.3229460158294657   0.9634637873769205   0.49703152004709966   0.13707247740226033   0.5685677129379152   0.836941647960681   0.5571619979252764   0.5981034971815041   0.3985578506112502   0.0725897164693207   0.5161054240968411   0.8963620333461885   0.2042038383748401   0.11984406339644002
0.46189137246009465   0.6555066192142189   0.011797688439479549   0.7494380907326773   0.5765745991980019   0.6465558148431099   0.20896616472498508   0.9262377988082239   0.3482858478849038   0.5884450496101218   0.8860201488955194   0.9627740114313034   0.8512543278378042   0.4513725722078614   0.31745243595760425   0.12583236347062235   0.29409232991252776   0.8532690750263573   0.918894585346354   0.05324264700130165   0.7779869058156866   0.9569070416801688   0.7146907469715139   0.9333985836048616   0.316095533355592   0.3014004224659499   0.7028930585320344   0.18396049287218436   0.73952093415759   0.65484460762284   0.4939268938070493   0.2577226940639604   0.3912350862726862   0.06639955801271832   0.6079067449115299   0.29494868263265706   0.539980758434882   0.6150269858048569   0.29045430895392566   0.16911631916203468   0.24588842852235432   0.7617579107784996   0.3715597236075716   0.11587367216073303   0.46790152270666774   0.8048508690983307   0.6568689766360577   0.1824750885558714   0.15180598935107575   0.5034504466323808   0.9539759181040233   0.9985145956836871   0.41228505519348574   0.8486058390095408   0.46004902429697403   0.7407919016197266   0.02104996892079951   0.7822062809968224   0.8521422793854441   0.4458432189870696   0.48106921048591744   0.16717929519196553   0.5616879704315184   0.2767268998250349
0.23518078196356312   0.405421384413466   0.19012824682394686   0.16085322766430185   0.7672792592568954   0.6005705153151352   0.5332592701878892   0.9783781391084304   0.6154732699058196   0.09712006868275438   0.5792833520838658   0.9798635434247434   0.20318821471233392   0.24851422967321363   0.11923432778689184   0.23907164180501675   0.18213824579153443   0.4663079486763912   0.26709204840144773   0.7932284228179471   0.7010690353056169   0.2991286534844257   0.7054040779699293   0.5165015229929123   0.46588825334205386   0.8937072690709598   0.5152758311459824   0.3556482953286104   0.6986089940851584   0.2931367537558245   0.9820165609580933   0.37727015622018   0.08313572417933882   0.1960166850730701   0.4027332088742274   0.3974066127954366   0.8799475094670048   0.9475024553998564   0.28349888108733556   0.15833497099041988   0.6978092636754705   0.48119450672346525   0.016406832685887846   0.3651065481724727   0.9967402283698535   0.1820658532390396   0.31100275471595856   0.8486050251795604   0.5308519750277997   0.28835858416807986   0.7957269235699761   0.49295672985094996   0.8322429809426412   0.9952218304122554   0.8137103626118829   0.11568657363076996   0.7491072567633024   0.7992051453391853   0.4109771537376555   0.7182799608353333   0.8691597472962975   0.8517026899393288   0.12747827265031986   0.5599449898449135
0.171350483620827   0.37050818321586354   0.11107143996443203   0.1948384416724408   0.17461025525097348   0.18844232997682395   0.8000686852484734   0.34623341649288036   0.6437582802231738   0.9000837458087441   0.00434176167849731   0.8532766866419305   0.8115152992805327   0.9048619153964886   0.19063139906661444   0.7375901130111605   0.06240804251723027   0.10565677005730341   0.779654245328959   0.019310152175827117   0.1932482952209328   0.2539540801179746   0.6521759726786391   0.4593651623309136   0.02189781160010579   0.8834458969021111   0.5411045327142071   0.2645267206584729   0.8472875563491323   0.6950035669252871   0.7410358474657336   0.9182933041655925   0.20352927612595847   0.794919821116543   0.7366940857872364   0.06501661752366204   0.3920139768454258   0.8900579057200544   0.5460626867206219   0.3274265045125016   0.32960593432819557   0.7844011356627509   0.7664084413916629   0.30811635233667445   0.13635763910726276   0.5304470555447763   0.11423246871302378   0.8487511900057608   0.11445982750715697   0.6470011586426653   0.5731279359988167   0.584224469347288   0.26717227115802467   0.9519975917173782   0.832092088533083   0.6659311651816955   0.0636429950320662   0.15707777060083514   0.09539800274584671   0.6009145476580334   0.6716290181866403   0.2670198648807808   0.5493353160252248   0.2734880431455319
0.3420230838584448   0.48261872921802984   0.7829268746335619   0.9653716908088574   0.20566544475118206   0.9521716736732535   0.6686944059205381   0.11662050080309658   0.09120561724402511   0.3051705150305883   0.09556646992172145   0.5323960314558086   0.8240333460860004   0.3531729233132101   0.2634743813886384   0.8664648662741131   0.7603903510539343   0.196095152712375   0.16807637864279168   0.26555031861607964   0.08876133286729385   0.9290752878315942   0.6187410626175669   0.9920622754705478   0.746738249008849   0.44645655861356437   0.835814187984005   0.026690584661690362   0.5410728042576669   0.4942848849403108   0.16711978206346684   0.9100700838585938   0.4498671870136418   0.18911436990972255   0.07155331214174539   0.3776740524027852   0.6258338409276414   0.8359414465965125   0.808078930753107   0.511209186128672   0.8654434898737072   0.6398462938841375   0.6400025521103153   0.24565886751259247   0.7766821570064133   0.7107710060525433   0.021261489492748423   0.2535965920420447   0.029943907997564315   0.2643144474389789   0.18544730150874347   0.22690600738035435   0.4888711037398974   0.770029562498668   0.018327519445276642   0.31683592352176054   0.039003916726255534   0.5809151925889455   0.9467742073035312   0.9391618711189753   0.41317007579861414   0.744973745992433   0.13869527655042427   0.42795268499030326
0.547726585924907   0.10512745210829563   0.498692724440109   0.18229381747771078   0.7710444289184937   0.3943564460557524   0.47743123494736056   0.9286972254356661   0.7411005209209293   0.13004199861677346   0.2919839334386171   0.7017912180553117   0.2522294171810319   0.36001243611810535   0.27365641399334045   0.3849552945335512   0.2132255004547764   0.7790972435291598   0.32688220668980916   0.44579342341457584   0.8000554246561623   0.034123497536726714   0.18818693013938492   0.017840738424272595   0.25232883873125533   0.9289960454284311   0.6894942056992759   0.8355469209465618   0.48128440981276166   0.5346395993726787   0.21206297075191538   0.9068496955108957   0.7401838888918324   0.4045976007559053   0.9200790373132983   0.20505847745558395   0.4879544717108004   0.04458516463779993   0.6464226233199578   0.8201031829220328   0.274728971256024   0.2654879211086401   0.31954041663014865   0.37430975950745693   0.4746735465998618   0.23136442357191342   0.13135348649076373   0.3564690210831843   0.22234470786860647   0.30236837814348233   0.4418592807914878   0.5209221001366225   0.7410602980558448   0.7677287787708036   0.22979631003957243   0.6140724046257268   0.0008764091640124068   0.3631311780148983   0.30971727272627414   0.40901392717014284   0.512921937453212   0.31854601337709837   0.6632946494063163   0.5889107442481101
0.2381929661971879   0.05305809226845827   0.3437542327761677   0.21460098474065317   0.7635194195973262   0.8216936686965448   0.21240074628540395   0.8581319636574689   0.5411747117287197   0.5193252905530625   0.7705414654939162   0.33720986352084636   0.8001144136728748   0.751596511782259   0.5407451554543438   0.7231374588951196   0.7992380045088625   0.3884653337673606   0.2310278827280696   0.3141235317249767   0.2863160670556505   0.06991932039026222   0.5677332333217533   0.7252127874768667   0.048123100858462595   0.01686122812180395   0.2239790005455856   0.5106118027362134   0.28460368126113644   0.1951675594252591   0.011578254260181628   0.6524798390787446   0.7434289695324168   0.6758422688721966   0.24103678876626547   0.31526997555789826   0.9433145558595419   0.9242457570899376   0.7002916333119217   0.5921325166627787   0.14407655135067943   0.535780423322577   0.4692637505838521   0.278008984937802   0.8577604842950289   0.46586110293231475   0.9015305172620989   0.5527961974609353   0.8096373834365663   0.44899987481051085   0.6775515167165133   0.042184394724721914   0.5250337021754299   0.25383231538525175   0.6659732624563316   0.38970455564597734   0.7816047326430131   0.5779900465130552   0.42493647369006615   0.07443458008807906   0.8382901767834712   0.6537442894231176   0.7246448403781445   0.48230206342530035
0.6942136254327917   0.11796386610054058   0.2553810897942923   0.20429307848749836   0.8364531411377628   0.6521027631682258   0.3538505725321935   0.651496881026563   0.026815757701196465   0.20310288835771498   0.6762990558156802   0.6093124863018411   0.5017820555257666   0.9492705729724632   0.010325793359348582   0.21960793065586376   0.7201773228827535   0.37128052645940807   0.5853893196692824   0.14517335056778471   0.8818871460992823   0.7175362370362904   0.860744479291138   0.6628712871424843   0.18767352066649062   0.5995723709357499   0.6053633894968456   0.458578208654986   0.3512203795287278   0.9474696077675241   0.25151281696465216   0.807081327628423   0.3244046218275314   0.7443667194098091   0.5752137611489719   0.19776884132658193   0.8226225663017648   0.7950961464373459   0.5648879677896234   0.9781609106707182   0.10244524341901125   0.4238156199779379   0.9794986481203409   0.8329875601029335   0.22055809731972892   0.7062793829416474   0.11875416882920298   0.17011627296044912   0.03288457665323829   0.1067070120058975   0.5133907793323573   0.7115380643054632   0.6816641971245104   0.1592374042383734   0.2618779623677052   0.9044567366770401   0.3572595752969791   0.41487068482856426   0.6866642012187333   0.7066878953504582   0.5346370089952144   0.6197745383912184   0.12177623342910995   0.72852698467974
0.4321917655762031   0.19595891841328053   0.14227758530876902   0.8955394245768065   0.2116336682564742   0.4896795354716331   0.023523416479566045   0.7254231516163574   0.1787490916032359   0.3829725234657357   0.5101326371472087   0.01388508731089426   0.49708489447872545   0.22373511922736225   0.24825467477950347   0.10942835063385414   0.13982531918174634   0.808864434398798   0.5615904735607702   0.40274045528339597   0.605188310186532   0.18908989600757958   0.4398142401316602   0.674213470603656   0.1729965446103289   0.993130977594299   0.2975366548228912   0.7786740460268494   0.9613628763538548   0.5034514421226659   0.27401323834332514   0.05325089441049207   0.7826137847506188   0.12047891865693025   0.7638806011961164   0.039365807099597805   0.2855288902718934   0.8967437994295681   0.515625926416613   0.9299374564657437   0.14570357109014703   0.08787936503077003   0.9540354528558428   0.5271970011823477   0.540515260903615   0.8987894690231905   0.5142212127241826   0.8529835305786917   0.36751871629328614   0.9056584914288913   0.21668455790129143   0.07430948455184226   0.40615583993943144   0.4022070493062255   0.9426713195579662   0.02105859014135019   0.6235420551888127   0.2817281306492952   0.17879071836184982   0.9816927830417523   0.3380131649169193   0.3849843312197272   0.6631647919452368   0.05175532657600872
0.19230959382677226   0.29710496618895715   0.709129339089394   0.524558325393661   0.6517943329231572   0.39831549716576675   0.1949081263652114   0.6715747948149693   0.28427561662987105   0.4926570057368754   0.97822356846392   0.597265310263127   0.8781197766904396   0.0904499564306499   0.0355522489059537   0.5762067201217769   0.25457772150162694   0.8087218257813547   0.8567615305441039   0.5945139370800244   0.9165645565847077   0.4237374945616275   0.19359673859886706   0.5427586105040157   0.7242549627579354   0.12663252837267033   0.48446739950947304   0.01820028511035473   0.0724606298347782   0.7283170312069036   0.28955927314426166   0.3466254902953854   0.7881850132049072   0.2356600254700282   0.31133570468034166   0.7493601800322583   0.9100652365144676   0.1452100690393783   0.27578345577438795   0.17315345991048153   0.6554875150128406   0.3364882432580236   0.4190219252302841   0.578639522830457   0.7389229584281329   0.9127507486963962   0.22542518663141703   0.0358809123264413   0.014667995670197534   0.7861182203237258   0.740957787121944   0.017680627216086566   0.9422073658354193   0.0578011891168222   0.4513985139776823   0.6710551369207012   0.15402235263051217   0.822141163646794   0.14006280929734066   0.9216949568884427   0.24395711611604465   0.6769310946074156   0.8642793535229527   0.7485414969779612
0.588469601103204   0.34044285134939206   0.4452574282926686   0.1699019741475042   0.8495466426750711   0.42769210265299595   0.21983224166125157   0.1340210618210629   0.8348786470048736   0.6415738823292702   0.47887445453930755   0.11634043460497634   0.8926712811694543   0.583772693212448   0.027475940561625226   0.4452852976842752   0.738648928538942   0.7616315295656539   0.8874131312642846   0.5235903407958324   0.4946918124228974   0.0847004349582383   0.02313377774133187   0.7750488438178712   0.9062222113196934   0.7442575836088462   0.5778763494486633   0.605146869670367   0.05667556864462228   0.3165654809558503   0.3580441077874117   0.4711258078493041   0.22179692163974873   0.6749915986265802   0.8791696532481041   0.35478537324432774   0.3291256404702945   0.0912189054141322   0.851693712686479   0.9095000755600525   0.5904767119313524   0.32958737584847825   0.9642805814221944   0.38590973476422014   0.09578489950845506   0.24488694089023993   0.9411468036808625   0.610860890946349   0.18956268818876168   0.5006293572813937   0.3632704542321992   0.00571402127598198   0.1328871195441394   0.18406387632554336   0.005226346444787505   0.534588213426678   0.9110901979043907   0.5090722776989632   0.12605669319668336   0.17980284018235018   0.5819645574340961   0.417853372284831   0.2743629805102044   0.27030276462229763
0.9914878455027437   0.08826599643635277   0.31008239908801005   0.8843930298580776   0.8957029459942887   0.8433790555461128   0.36893559540714754   0.27353213891172856   0.706140257805527   0.3427496982647192   0.005665141174948348   0.2678181176357466   0.5732531382613876   0.1586858219391758   0.0004387947301608421   0.7332299042090686   0.6621629403569969   0.6496135442402126   0.8743821015334775   0.5534270640267185   0.08019838292290071   0.23176017195538157   0.600019121023273   0.28312429940442085   0.08871053742015698   0.1434941755190288   0.289936721935263   0.39873126954634336   0.19300759142586832   0.30011511997291596   0.9210011265281154   0.12519913063461482   0.48686733362034135   0.9573654217081968   0.9153359853531671   0.8573810129988683   0.9136141953589537   0.798679599769021   0.9148971906230062   0.1241511087897996   0.25145125500195686   0.1490660555288084   0.04051508908952875   0.5707240447630811   0.17125287207905615   0.9173058835734268   0.4404959680662557   0.28759974535866023   0.08254233465889917   0.773811708054398   0.1505592461309927   0.8888684758123169   0.8895347432330308   0.4736965880814821   0.22955811960287728   0.7636693451777021   0.40266740961268954   0.5163311663732852   0.3142221342497102   0.9062883321788339   0.48905321425373577   0.7176515666042643   0.39932494362670395   0.7821372233890342
0.2376019592517789   0.568585511075456   0.35880985453717523   0.2114131786259531   0.06634908717272275   0.6512796275020291   0.9183138864709195   0.9238134332672928   0.9838067525138235   0.877467919447631   0.7677546403399268   0.034944957454975965   0.09427200928079274   0.403771331366149   0.5381965207370496   0.27127561227727387   0.6916045996681032   0.8874401649928637   0.22397438648733936   0.36498728009844006   0.20255138541436746   0.16978859838859942   0.8246494428606354   0.5828500567094058   0.9649494261625885   0.6012030873131435   0.4658395883234602   0.3714368780834527   0.8986003389898658   0.9499234598111144   0.5475257018525407   0.44762344481615984   0.9147935864760423   0.07245554036348334   0.7797710615126139   0.4126784873611839   0.8205215771952494   0.6686842089973344   0.24157454077556428   0.14140287508391   0.12891697752714626   0.7812440440044707   0.01760015428822492   0.77641559498547   0.9263655921127788   0.6114554456158712   0.19295071142758952   0.19356553827606413   0.9614161659501903   0.010252358302727697   0.7271111231041293   0.8221286601926114   0.06281582696032446   0.06032889849161328   0.17958542125158866   0.37450521537645154   0.14802224048428225   0.9878733581281299   0.39981435973897483   0.9618267280152677   0.32750066328903277   0.3191891491307956   0.15823981896341052   0.8204238529313577
0.1985836857618865   0.537945105126325   0.14063966467518563   0.04400825794588768   0.2722180936491077   0.9264896595104538   0.947688953247596   0.8504427196698235   0.31080192769891746   0.9162373012077261   0.22057783014346677   0.028314059477212154   0.24798610073859298   0.8559084027161128   0.04099240889187812   0.6538088441007606   0.09996386025431073   0.8680350445879829   0.6411780491529033   0.691982116085493   0.772463196965278   0.5488458954571873   0.4829382301894928   0.8715582631541353   0.5738795112033914   0.010900790330862288   0.34229856551430715   0.8275500052082476   0.3016614175542837   0.08441113082040852   0.39460961226671104   0.9771072855384241   0.9908594898553663   0.16817382961268243   0.17403178212324427   0.9487932260612119   0.7428733891167734   0.31226542689656966   0.13303937323136614   0.2949843819604513   0.6429095288624627   0.4442303823085868   0.49186132407846284   0.6030022658749583   0.8704463318971847   0.8953844868513995   0.008923093888970076   0.731444002720823   0.2965668206937932   0.8844836965205373   0.6666245283746629   0.9038939975125754   0.9949054031395095   0.8000725657001287   0.27201491610795187   0.9267867119741513   0.004045913284143166   0.6318987360874463   0.09798313398470761   0.9779934859129394   0.26117252416736986   0.3196333091908766   0.9649437607533414   0.6830091039524882
0.6182629953049072   0.8754029268822898   0.4730824366748786   0.08000683807752978   0.7478166634077226   0.9800184400308903   0.46415934278590854   0.34856283535670674   0.45124984271392937   0.09553474351035311   0.7975348144112456   0.4446688378441313   0.4563444395744199   0.2954621778102244   0.5255198983032937   0.51788212586998   0.4522985262902767   0.6635634417227781   0.4275367643185861   0.5398886399570405   0.19112600212290687   0.34393013253190147   0.4625930035652447   0.8568795360045524   0.5728630068179996   0.46852720564961164   0.9895105668903661   0.7768726979270226   0.825046343410277   0.4885087656187213   0.5253512241044576   0.4283098625703159   0.37379650069634773   0.3929740221083682   0.7278164096932119   0.9836410247261845   0.9174520611219279   0.09751184429814377   0.2022965113899182   0.4657588988562046   0.46515353483165117   0.43394840257536565   0.7747597470713321   0.925870258899164   0.2740275327087443   0.09001827004346416   0.31216674350608736   0.06899072289461161   0.7011645258907446   0.6214910643938525   0.3226561766157213   0.292118024967589   0.8761181824804676   0.13298229877513124   0.7973049525112638   0.8638081623972731   0.5023216817841198   0.740008276666763   0.06948854281805186   0.8801671376710886   0.584869620662192   0.6424964323686193   0.8671920314281336   0.41440823881488403
0.11971608583054079   0.20854802979325363   0.0924322843568016   0.48853797991572   0.8456885531217965   0.11852975974978947   0.7802655408507142   0.4195472570211084   0.14452402723105187   0.4970386953559369   0.4576093642349929   0.1274292320535194   0.2684058447505843   0.3640563965808057   0.6603044117237291   0.26362106965624627   0.7660841629664645   0.6240481199140426   0.5908158689056773   0.38345393198515765   0.18121454230427256   0.9815516875454234   0.7236238374775436   0.9690456931702737   0.061498456473731776   0.7730036577521697   0.6311915531207419   0.48050771325455366   0.21580990335193526   0.6544738980023803   0.8509260122700277   0.06096045623344527   0.0712858761208834   0.15743520264644337   0.39331664803503485   0.9335312241799258   0.8028800313702991   0.7933788060656376   0.7330122363113057   0.6699101545236796   0.03679586840383456   0.169330686151595   0.1421963674056285   0.28645622253852193   0.855581326099562   0.18777899860617162   0.4185725299280849   0.3174105293682483   0.7940828696258302   0.41477534085400186   0.7873809768073429   0.8369028161136947   0.5782729662738949   0.7603014428516216   0.9364549645373151   0.7759423598802494   0.5069870901530116   0.6028662402051782   0.5431383165022803   0.8424111357003234   0.7041070587827125   0.8094874341395405   0.8101260801909745   0.17250098117664384
0.6673111903788779   0.6401567479879455   0.6679297127853461   0.8860447586381219   0.8117298642793159   0.45237774938177394   0.24935718285726116   0.5686342292698736   0.017646994653485702   0.03760240852777208   0.4619762060499183   0.731731413156179   0.4393740283795908   0.27730096567615053   0.5255212415126032   0.9557890532759296   0.9323869382265793   0.6744347254709724   0.9823829250103229   0.11337791757560609   0.2282798794438667   0.8649472913314318   0.1722568448193483   0.9408769363989622   0.5609686890649888   0.22479054334348625   0.5043271320340023   0.054832177760840345   0.7492388247856728   0.7724127939617124   0.25496994917674104   0.48619794849096676   0.7315918301321872   0.7348103854339403   0.7929937431268228   0.7544665353347878   0.29221780175259643   0.4575094197577897   0.26747250161421965   0.7986774820588582   0.35983086352601723   0.7830746942868174   0.28508957660389683   0.6852995644832521   0.1315509840821505   0.9181274029553855   0.11283273178454853   0.7444226280842899   0.5705822950171617   0.6933368596118993   0.6085055997505463   0.6895904503234496   0.8213434702314888   0.920924065650187   0.3535356505738052   0.20339250183248284   0.08975164009930163   0.18611368021624675   0.5605419074469824   0.448925966497695   0.7975338383467052   0.728604260458457   0.29306940583276275   0.6502484844388368
0.437702974820688   0.9455295661716396   0.007979829228865924   0.9649489199555846   0.3061519907385375   0.02740216321625408   0.8951470974443174   0.22052629187129466   0.7355696957213758   0.33406530360435477   0.2866414976937711   0.5309358415478451   0.914226225489887   0.4131412379541678   0.9331058471199659   0.32754333971536226   0.8244745853905854   0.22702755773792102   0.37256393967298346   0.8786173732176672   0.02694074704388015   0.498423297279464   0.0794945338402207   0.22836888877883046   0.5892377722231922   0.5528937311078244   0.07151470461135478   0.26341996882324586   0.2830857814846547   0.5254915678915703   0.1763676071670374   0.042893676951951204   0.5475160857632789   0.1914262642872155   0.8897261094732662   0.5119578354041061   0.633289860273392   0.7782850263330477   0.9566202623533004   0.18441449568874388   0.8088152748828066   0.5512574685951267   0.5840563226803169   0.30579712247107665   0.7818745278389264   0.05283417131566269   0.5045617888400963   0.07742823369224619   0.19263675561573423   0.49994044020783834   0.43304708422874144   0.8140082648690004   0.9095509741310795   0.9744488723162681   0.2566794770617041   0.7711145879170491   0.3620348883678007   0.7830226080290525   0.3669533675884378   0.259156752512943   0.7287450280944088   0.004737581696004856   0.4103331052351374   0.07474225682419912
0.9199297532116022   0.45348011310087816   0.8262767825548204   0.7689451343531225   0.13805522537267576   0.40064594178521545   0.32171499371472423   0.6915169006608762   0.9454184697569415   0.9007055015773772   0.8886679094859827   0.877508635791876   0.03586749562586196   0.9262566292611091   0.6319884324242787   0.10639404787482683   0.6738326072580613   0.14323402123205647   0.26503506483584094   0.8472372953618839   0.9450875791636526   0.13849643953605162   0.8547019596007035   0.7724950385376848   0.0251578259520504   0.6850163264351735   0.028425177045883102   0.00354990418456226   0.8871026005793746   0.284370384649958   0.7067101833311589   0.312033003523686   0.9416841308224331   0.38366488307258084   0.8180422738451761   0.43452436773181   0.9058166351965712   0.45740825381147177   0.18605384142089745   0.3281303198569832   0.23198402793850986   0.3141742325794153   0.9210187765850565   0.48089302449509935   0.28689644877485726   0.17567779304336367   0.06631681698435299   0.7083979859574147   0.2617386228228069   0.4906614666081902   0.03789163993846989   0.7048480817728524   0.37463602224343223   0.20629108195823223   0.33118145660731096   0.3928150782491664   0.4329518914209991   0.8226261988856514   0.5131391827621349   0.9582907105173564   0.5271352562244279   0.3652179450741796   0.3270853413412374   0.6301603906603731
0.2951512282859181   0.05104371249476429   0.40606656475618086   0.14926736616527378   0.008254779511060815   0.8753659194514006   0.33974974777182787   0.4408693802078591   0.7465161566882539   0.3847044528432104   0.301858107833358   0.7360212984350067   0.37188013444482165   0.1784133708849782   0.970676651226047   0.3432062201858403   0.9389282430238226   0.3557871719993268   0.45753746846391213   0.3849155096684839   0.4117929867993946   0.9905692269251472   0.13045212712267476   0.7547551190081108   0.1166417585134765   0.9395255144303829   0.7243855623664939   0.605487752842837   0.10838697900241567   0.06415959497898228   0.384635814594666   0.1646183726349779   0.36187082231416173   0.6794551421357719   0.08277770676130804   0.4285970741999712   0.9899906878693401   0.5010417712507937   0.11210105553526103   0.08539085401413087   0.051062444845517516   0.14525459925146691   0.6545635870713489   0.700475344345647   0.6392694580461229   0.1546853723263197   0.5241114599486741   0.9457202253375361   0.5226276995326464   0.2151598578959368   0.7997258975821803   0.3402324724946991   0.41424072053023075   0.1510002629169545   0.41509008298751426   0.17561409985972123   0.05236989821606901   0.4715451207811826   0.33231237622620624   0.74701702565975   0.06237921034672894   0.970503349530389   0.22021132069094518   0.6616261716456192
0.011316765501211428   0.825248750278922   0.5656477336195963   0.9611508272999723   0.3720473074550885   0.6705633779526023   0.041536273670922136   0.015430601962436155   0.8494196079224421   0.4554035200566655   0.24181037608874187   0.675198129467737   0.43517888739221133   0.304403257139711   0.8267202931012276   0.4995840296080158   0.3828089891761423   0.8328581363585283   0.4944079168750214   0.7525670039482657   0.32042977882941337   0.8623547868281395   0.2741965961840762   0.09094083230264652   0.30911301332820196   0.03710603654921745   0.7085488625644799   0.12979000500267424   0.9370657058731134   0.36654265859661517   0.6670125888935579   0.11435940304023808   0.08764609795067135   0.9111391385399497   0.42520221280481596   0.43916127357250107   0.65246721055846   0.6067358814002386   0.5984819197035883   0.9395772439644853   0.2696582213823177   0.7738777450417103   0.1040740028285669   0.18701024001621952   0.9492284425529044   0.9115229582135708   0.8298774066444906   0.096069407713573   0.6401154292247024   0.8744169216643534   0.1213285440800107   0.9662794027108987   0.703049723351589   0.5078742630677382   0.4543159551864529   0.8519199996706607   0.6154036254009176   0.5967351245277885   0.029113742381636942   0.4127587260981596   0.9629364148424576   0.9899992431275499   0.4306318226780486   0.4731814821336744
0.6932781934601399   0.21612149808583966   0.32655781984948173   0.28617124211745487   0.7440497509072355   0.30459853987226887   0.49668041320499107   0.19010183440388184   0.1039343216825331   0.4301816182079155   0.37535186912498036   0.22382243169298308   0.40088459833094414   0.9223073551401773   0.9210359139385275   0.3719024320223224   0.7854809729300265   0.3255722306123887   0.8919221715568906   0.9591437059241628   0.8225445580875689   0.33557298748483877   0.4612903488788419   0.48596222379048837   0.12926636462742905   0.11945148939899912   0.1347325290293602   0.19979098167303355   0.3852166137201935   0.8148529495267303   0.6380521158243692   0.00968914726915169   0.2812822920376604   0.38467133131881476   0.26270024669938874   0.7858667155761686   0.8803976937067163   0.46236397617863745   0.3416643327608612   0.4139642835538462   0.09491672077668979   0.13679174556624873   0.4497421612039707   0.4548205776296834   0.2723721626891209   0.80121875808141   0.9884518123251288   0.968858353839195   0.14310579806169185   0.6817672686824108   0.8537192832957685   0.7690673721661615   0.7578891843414983   0.8669143191556806   0.21566716747139947   0.7593782248970098   0.4766068923038379   0.4822429878368658   0.9529669207720107   0.9735115093208412   0.5962091985971216   0.019879011658228345   0.6113025880111495   0.559547225766995
0.5012924778204318   0.8830872660919796   0.1615604268071788   0.10472664813731157   0.22892031513131095   0.08186850801056965   0.17310861448205006   0.13586829429811653   0.08581451706961908   0.40010123932815883   0.3193893311862815   0.36680092213195503   0.32792533272812074   0.5331869201724783   0.10372216371488202   0.6074226972349452   0.8513184404242828   0.05094393233561244   0.1507552429428713   0.6339111879141041   0.25510924182716116   0.03106492067738409   0.5394526549317218   0.07436396214710905   0.7538167640067294   0.1479776545854045   0.377892228124543   0.9696373140097975   0.5248964488754184   0.06610914657483484   0.20478361364249292   0.8337690197116809   0.43908193180579935   0.666007907246676   0.8853942824562114   0.4669680975797259   0.1111565990776786   0.1328209870741978   0.7816721187413295   0.8595454003447807   0.25983815865339577   0.08187705473858534   0.6309168757984581   0.22563421243067658   0.004728916826234606   0.05081213406120125   0.09146422086673635   0.15127025028356753   0.25091215281950524   0.9028344794757968   0.7135719927421934   0.18163293627377006   0.7260157039440869   0.836725332900962   0.5087883790997004   0.3478639165620891   0.2869337721382875   0.1707174256542859   0.623394096643489   0.8808958189823632   0.17577717306060892   0.03789643858008813   0.8417219779021595   0.02135041863758259
0.9159390144072131   0.9560193838415028   0.21080510210370143   0.795716206206906   0.9112100975809785   0.9052072497803015   0.1193408812369651   0.6444459559233384   0.6602979447614733   0.0023727703045047744   0.4057688884947717   0.46281301964956845   0.9342822408173864   0.16564743740354285   0.8969805093950712   0.11494910308747931   0.6473484686790989   0.994930011749257   0.2735864127515823   0.23405328410511608   0.47157129561849   0.9570335731691688   0.4318644348494227   0.2127028654675335   0.5556322812112768   0.0010141893276660397   0.2210593327457213   0.4169866592606275   0.6444221836302984   0.09580693954736451   0.10171845150875618   0.772540703337289   0.984124238868825   0.09343416924285973   0.6959495630139845   0.3097276836877206   0.04984199805143861   0.9277867318393169   0.7989690536189131   0.19477858060024128   0.40249352937233973   0.9328567200900599   0.5253826408673309   0.9607252964951252   0.9309222337538497   0.9758231469208911   0.09351820601790817   0.7480224310275917   0.37528995254257286   0.9748089575932251   0.8724588732721869   0.3310357717669642   0.7308677689122746   0.8790020180458605   0.7707404217634307   0.5584950684296752   0.7467435300434495   0.7855678488030008   0.07479085874944626   0.24876738474195462   0.696901531992011   0.857781116963684   0.27582180513053306   0.05398880414171332
0.29440800261967126   0.924924396873624   0.7504391642632022   0.09326350764658814   0.3634857688658215   0.9491012499527329   0.6569209582452941   0.34524107661899645   0.9881958163232486   0.9742922923595079   0.7844620849731071   0.014205304852032228   0.25732804741097404   0.09529027431364731   0.01372166320967642   0.45571023642235703   0.5105845173675245   0.3097224255106465   0.9389308044602301   0.20694285168040244   0.8136829853755135   0.4519413085469625   0.6631089993296971   0.1529540475386891   0.5192749827558423   0.5270169116733385   0.9126698350664949   0.05969053989210098   0.15578921389002082   0.5779156617206056   0.25574887682120084   0.7144494632731045   0.1675933975667722   0.6036233693610977   0.47128679184809374   0.7002441584210723   0.9102653501557981   0.5083330950474504   0.4575651286384173   0.24453392199871526   0.39968083278827365   0.19861066953680392   0.5186343241781871   0.03759107031831284   0.5859978474127601   0.7466693609898414   0.8555253248484901   0.8846370227796237   0.06672286465691776   0.21965244931650288   0.9428554897819952   0.8249464828875228   0.9109336507668969   0.6417367875958973   0.6871066129607943   0.11049701961441823   0.7433402532001248   0.03811341823479959   0.21581982111270057   0.4102528611933459   0.8330749030443266   0.5297803231873492   0.7582546924742832   0.16571893919463063
0.4333940702560529   0.3311696536505453   0.23962036829609612   0.1281278688763178   0.8473962228432929   0.5845002926607039   0.3840950434476061   0.24349084609669405   0.7806733581863751   0.364847843344201   0.4412395536656109   0.4185443632091713   0.8697397074194781   0.7231110557483037   0.7541329407048166   0.3080473435947531   0.1263994542193534   0.6849976375135041   0.538313119592116   0.8977944824014071   0.29332455117502676   0.1552173143261549   0.7800584271178328   0.7320755432067765   0.8599304809189738   0.8240476606756096   0.5404380588217367   0.6039476743304587   0.012534258075680975   0.23954736801490575   0.15634301537413056   0.3604568282337647   0.2318608998893059   0.8746995246707048   0.7151034617085197   0.9419124650245934   0.36212119246982777   0.15158846892240105   0.9609705210037031   0.6338651214298403   0.23572173825047438   0.46659083140889696   0.42265740141158703   0.7360706390284331   0.9423971870754476   0.311373517082742   0.6425989742937542   0.003995095821656576   0.08246670615647377   0.48732585640713244   0.10216091547201765   0.4000474214911978   0.0699324480807928   0.24777848839222666   0.9458179000978871   0.03959059325743317   0.8380715481914869   0.3730789637215219   0.23071443838936742   0.0976781282328398   0.47595035572165917   0.22149049479912086   0.26974391738566433   0.46381300680299953
0.24022861747118476   0.7548996633902239   0.8470865159740774   0.7277423677745665   0.2978314303957372   0.44352614630748183   0.20448754168032302   0.7237472719529099   0.21536472423926342   0.9562002899003494   0.10232662620830538   0.323699850461712   0.14543227615847062   0.7084218015081227   0.1565087261104183   0.2841092572042788   0.3073607279669837   0.33534283778660084   0.9257942877210509   0.18643112897143901   0.8314103722453245   0.11385234298748   0.6560503703353865   0.7226181221684395   0.5911817547741398   0.35895267959725613   0.8089638543613092   0.9948757543938731   0.2933503243784026   0.9154265332897743   0.6044763126809862   0.2711284824409632   0.07798560013913919   0.9592262433894249   0.5021496864726808   0.9474286319792512   0.9325533239806686   0.2508044418813021   0.3456409603622625   0.6633193747749724   0.6251925960136848   0.9154616040947012   0.4198466726412116   0.47688824580353334   0.7937822237683603   0.8016092611072212   0.7637963023058251   0.7542701236350938   0.20260046899422052   0.4426565815099651   0.9548324479445158   0.7593943692412208   0.9092501446158179   0.5272300482201908   0.35035613526352966   0.48826588680025756   0.8312645444766787   0.568003804830766   0.8482064487908488   0.5408372548210064   0.8987112204960102   0.31719936294946394   0.5025654884285863   0.8775178800460339
0.2735186244823253   0.4017377588547627   0.0827188157873747   0.4006296342425006   0.479736400713965   0.6001284977475415   0.3189225134815496   0.6463595106074067   0.2771359317197445   0.1574719162375764   0.3640900655370337   0.886965141366186   0.36788578710392655   0.6302418680173856   0.01373393027350404   0.39869925456592836   0.5366212426272479   0.06223806318661955   0.1655274814826552   0.8578619997449219   0.6379100221312377   0.7450387002371556   0.6629619930540689   0.980344119698888   0.36439139764891243   0.3433009413823929   0.5802431772666942   0.5797144854563874   0.8846549969349474   0.7431724436348514   0.26132066378514457   0.9333549748489807   0.6075190652152029   0.585700527397275   0.8972305982481108   0.04638983348279473   0.2396332781112764   0.9554586593798895   0.8834966679746068   0.6476905789168664   0.7030120354840286   0.8932205961932699   0.7179691864919516   0.7898285791719444   0.06510201335279088   0.14818189595611428   0.05500719343788277   0.8094844594730564   0.7007106157038785   0.8048809545737213   0.47476401617118863   0.229769974016669   0.8160556187689311   0.061708510938869976   0.21344335238604406   0.2964149991676883   0.20853655355372808   0.47600798354159496   0.3162127541379332   0.2500251656848936   0.9689032754424517   0.5205493241617055   0.4327160861633264   0.6023345867680272
0.2658912399584231   0.6273287279684356   0.7147468996713748   0.8125060075960828   0.20078922660563223   0.47914683201232133   0.659739706233492   0.0030215481230264248   0.5000786109017538   0.6742658774386   0.1849756900623034   0.7732515741063575   0.6840229921328227   0.61255736649973   0.9715323376762593   0.4768365749386691   0.4754864385790946   0.136549382958135   0.6553195835383262   0.2268114092537755   0.506583163136643   0.6160000587964295   0.22260349737499974   0.6244768224857483   0.24069192317821983   0.9886713308279939   0.507856597703625   0.8119708148896655   0.039902696572587604   0.5095244988156725   0.8481168914701329   0.808949266766639   0.5398240856708338   0.8352586213770725   0.6631412014078295   0.035697692660281596   0.8558010935380111   0.22270125487734252   0.6916088637315702   0.5588611177216125   0.3803146549589166   0.08615187191920749   0.03628928019324403   0.332049708467837   0.8737314918222736   0.470151813122778   0.8136857828182443   0.7075728859820888   0.6330395686440539   0.48148048229478413   0.3058291851146193   0.8956020710924233   0.5931368720714663   0.9719559834791116   0.45771229364448635   0.08665280432578427   0.05331278640063235   0.13669736210203912   0.7945710922366568   0.05095511166550268   0.19751169286262119   0.9139961072246966   0.10296222850508664   0.4920939939438902
0.8171970379037046   0.8278442353054891   0.06667294831184262   0.16004428547605315   0.943465546081431   0.3576924221827111   0.25298716549359834   0.4524713994939644   0.31042597743737715   0.876211939887927   0.947157980378979   0.5568693284015411   0.717289105365911   0.9042559564088153   0.4894456867344926   0.4702165240757568   0.6639763189652786   0.7675585943067762   0.6948745944978358   0.41926141241025416   0.46646462610265743   0.8535624870820796   0.5919123659927492   0.927167418466364   0.6492675881989528   0.02571825177659052   0.5252394176809065   0.7671231329903109   0.7058020421175218   0.6680258295938795   0.2722522521873082   0.3146517334963464   0.39537606468014463   0.7918138897059525   0.3250942718083292   0.7577824050948053   0.6780869593142337   0.8875579332971372   0.8356485850738365   0.28756588101904845   0.014110640348955076   0.11999933899036096   0.14077399057600076   0.8683044686087943   0.5476460142462977   0.26643685190828137   0.5488616245832516   0.9411370501424303   0.8983784260473449   0.24071860013169083   0.023622206902345056   0.1740139171521195   0.19257638392982301   0.5726927705378114   0.7513699547150369   0.8593621836557731   0.7972003192496784   0.780878880831859   0.42627568290670764   0.10157977856096778   0.11911335993544468   0.8933209475347218   0.590627097832871   0.8140138975419193
0.10500271958648962   0.7733216085443608   0.4498531072568703   0.9457094289331249   0.557356705340192   0.5068847566360795   0.9009914826736187   0.004572378790694648   0.6589782792928471   0.26616615650438863   0.8773692757712737   0.8305584616385752   0.4664018953630241   0.6934733859665773   0.1259993210562368   0.9711962779828021   0.6692015761133457   0.9125945051347183   0.6997236381495292   0.8696164994218343   0.550088216177901   0.019273557599996535   0.10909654031665811   0.055602601879914976   0.44508549659141144   0.24595194905563572   0.6592434330597878   0.10989317294678999   0.8877287912512195   0.7390671924195563   0.7582519503861691   0.10532079415609534   0.22875051195837234   0.47290103591516763   0.8808826746148954   0.2747623325175202   0.7623486165953482   0.7794276499485904   0.7548833535586587   0.30356605453471813   0.09314704048200254   0.8668331448138721   0.05515971540912952   0.43394955511288386   0.5430588243041015   0.8475595872138756   0.9460631750924714   0.3783469532329689   0.09797332771269006   0.6016076381582398   0.2868197420326836   0.2684537802861789   0.2102445364614706   0.8625404457386836   0.5285677916465145   0.16313298613008356   0.9814940245030982   0.3896394098235159   0.647685117031619   0.8883706536125634   0.21914540790774997   0.6102117598749255   0.8928017634729604   0.5848045990778452
0.12599836742574744   0.7433786150610534   0.8376420480638308   0.15085504396496133   0.582939543121646   0.8958190278471778   0.8915788729713594   0.7725080907319924   0.4849662154089559   0.29421138968893795   0.6047591309386757   0.5040543104458135   0.27472167894748534   0.43167094395025435   0.07619133929216129   0.34092132431572997   0.2932276544443871   0.04203153412673843   0.4285062222605423   0.4525506707031666   0.07408224653663711   0.43181977425181295   0.535704458787582   0.8677460716253215   0.9480838791108896   0.6884411591907595   0.6980624107237512   0.7168910276603601   0.36514433598924373   0.7926221313435817   0.8064835377523918   0.9443829369283677   0.8801781205802878   0.49841074165464383   0.20172440681371603   0.44032862648255416   0.6054564416328024   0.06673979770438948   0.12553306752155474   0.09940730216682415   0.3122287871884154   0.024708263577651057   0.6970268452610124   0.6468566314636576   0.2381465406517783   0.5928884893258382   0.16132238647343047   0.7791105598383361   0.2900626615408886   0.9044473301350786   0.4632599757496793   0.062219532177976   0.9249183255516449   0.1118251987914968   0.6567764379972875   0.11783659524960834   0.0447402049713571   0.6134144571368529   0.45505203118357146   0.6775079687670542   0.4392837633385546   0.5466746594324635   0.3295189636620167   0.5781006666002301
0.12705497615013922   0.5219663958548124   0.6324921184010043   0.9312440351365725   0.888908435498361   0.9290779065289743   0.4711697319275738   0.1521334752982364   0.5988457739574723   0.02463057639389572   0.007909756177894505   0.0899139431202604   0.6739274484058274   0.9128053776023989   0.351133318180607   0.972077347870652   0.6291872434344703   0.29939092046554594   0.8960812869970356   0.2945693791035979   0.1899034800959157   0.7527162610330824   0.5665623233350189   0.7164687125033679   0.06284850394577648   0.23074986517827006   0.9340702049340146   0.7852246773667954   0.17394006844741555   0.30167195864929575   0.46290047300644077   0.633091202068559   0.5750942944899432   0.27704138225540004   0.45499071682854625   0.5431772589482985   0.9011668460841158   0.36423600465300116   0.10385739864793923   0.5710999110776465   0.2719796026496455   0.06484508418745517   0.20777611165090368   0.27653053197404864   0.08207612255372976   0.3121288231543727   0.6412137883158848   0.5600618194706808   0.019227618607953276   0.08137895797610264   0.7071435833818703   0.7748371421038854   0.8452875501605377   0.7797069993268069   0.24424311037542953   0.14174594003532653   0.2701932556705945   0.5026656170714068   0.7892523935468833   0.598568681087028   0.3690264095864787   0.1384296124184057   0.6853949948989441   0.02746877000938154
0.09704680693683325   0.07358452823095052   0.47761888324804036   0.7509382380353329   0.014970684383103483   0.7614557050765778   0.8364050949321555   0.19087641856465212   0.9957430657751503   0.6800767471004752   0.1292615115502852   0.41603927646076666   0.15045551561461248   0.9003697477736683   0.8850184011748556   0.2742933364254401   0.880262259944018   0.39770413070226146   0.09576600762797237   0.6757246553384121   0.5112358503575393   0.2592745182838558   0.4103710127290283   0.6482558853290306   0.414189043420706   0.18568999005290526   0.932752129480988   0.8973176472936977   0.3992183590376025   0.4242342849763274   0.09634703454883245   0.7064412287290455   0.4034752932624523   0.7441575378758523   0.9670855229985472   0.29040195226827886   0.25301977764783984   0.843787790102184   0.08206712182369158   0.016108615842838733   0.3727575177038219   0.4460836593999225   0.9863011141957192   0.34038396050442665   0.8615216673462827   0.18680914111606672   0.5759301014666909   0.6921280751753961   0.4473326239255766   0.0011191510631614633   0.6431779719857029   0.7948104278816984   0.04811426488797409   0.576884866086834   0.5468309374368705   0.08836919915265296   0.6446389716255218   0.8327273282109817   0.5797454144383233   0.7979672468843741   0.3916191939776819   0.9889395381087978   0.49767829261463165   0.7818586310415354
0.01886167627386006   0.5428558787088753   0.5113771784189125   0.44147467053710876   0.15734000892757743   0.3560467375928086   0.9354470769522216   0.7493465953617127   0.7100073850020008   0.3549275865296471   0.29226910496651864   0.9545361674800142   0.6618931201140268   0.7780427204428131   0.7454381675296482   0.8661669683273613   0.017254148488504976   0.9453153922318314   0.16569275309132495   0.06819972144298715   0.6256349545108231   0.9563758541230335   0.6680144604766933   0.2863410904014518   0.606773278236963   0.4135199754141582   0.15663728205778085   0.8448664198643431   0.44943326930938554   0.057473237821349624   0.22119020510555926   0.09551982450263037   0.7394258843073848   0.7025456512917025   0.9289211001390406   0.14098365702261617   0.07753276419335796   0.9245029308488893   0.18348293260939244   0.27481668869525494   0.06027861570485299   0.9791875386170581   0.017790179518067495   0.20661696725226777   0.4346436611940299   0.022811684494024514   0.3497757190413742   0.920275876850816   0.8278703829570669   0.6092917090798663   0.19313843698359337   0.07540945698647296   0.3784371136476814   0.5518184712585167   0.9719482318780341   0.9798896324838426   0.6390112293402967   0.8492728199668141   0.043027131738993474   0.8389059754612265   0.5614784651469388   0.9247698891179248   0.859544199129601   0.5640892867659715
0.5011998494420857   0.9455823505008667   0.8417540196115335   0.35747231951370373   0.06655618824805581   0.9227706660068422   0.49197830057015934   0.43719644266288776   0.23868580529098885   0.3134789569269759   0.298839863586566   0.36178698567641476   0.8602486916433074   0.7616604856684592   0.32689163170853186   0.3818973531925722   0.22123746230301072   0.9123876657016451   0.28386449996953844   0.5429913777313458   0.659758997156072   0.9876177765837203   0.4243203008399374   0.9789020909653743   0.15855914771398621   0.042035426082853544   0.5825662812284038   0.6214297714516706   0.0920029594659304   0.1192647600760113   0.09058798065824451   0.1842333287887828   0.8533171541749416   0.8057858031490354   0.7917481170716786   0.822446343112368   0.9930684625316342   0.0441253174805761   0.46485648536314667   0.44054898991979585   0.7718310002286234   0.13173765177893101   0.18099198539360825   0.8975576121884501   0.11207200307255143   0.14411987519521072   0.7566716845536708   0.9186555212230758   0.9535128553585652   0.10208444911235717   0.174105403325267   0.29722574977140526   0.8615098958926348   0.9828196890363459   0.08351742266702249   0.11299242098262248   0.008192741717693276   0.1770338858873105   0.291769305595344   0.29054607787025444   0.015124279186059164   0.1329085684067344   0.8269128202321973   0.8499970879504586
0.24329327895743577   0.0011709166278033852   0.6459208348385891   0.9524394757620086   0.13122127588488436   0.8570510414325927   0.8892491502849182   0.03378395453893278   0.17770842052631913   0.7549665923202356   0.7151437469596512   0.7365582047675275   0.3161985246336843   0.7721469032838897   0.6316263242926287   0.623565783784905   0.308005782915991   0.5951130173965792   0.33985701869728474   0.3330197059146506   0.2928815037299319   0.46220444898984475   0.5129441984650874   0.48302261796419194   0.0495882247724961   0.46103353236204137   0.8670233636264985   0.5305831422021834   0.9183669488876117   0.6039824909294487   0.9777742133415802   0.4967991876632506   0.7406585283612926   0.8490158986092132   0.26263046638192905   0.7602409828957231   0.42446000372760834   0.07686899532532356   0.6310041420893003   0.13667519911081805   0.11645422081161727   0.4817559779287444   0.2911471233920156   0.8036554931961675   0.8235727170816854   0.019551528938899658   0.7782029249269281   0.3206328752319755   0.7739844923091893   0.5585179965768583   0.9111795613004298   0.7900497330297921   0.8556175434215776   0.9545355056474096   0.9334053479588496   0.29325054536654155   0.11495901506028493   0.10551960703819639   0.6707748815769204   0.5330095624708184   0.6904990113326767   0.02865061171287284   0.039770739487620166   0.3963343633600004
0.5740447905210594   0.5468946337841284   0.7486236160956046   0.5926788701638329   0.7504720734393739   0.5273431048452287   0.9704206911686765   0.27204599493185744   0.9764875811301846   0.9688251082683704   0.059241129868246714   0.48199626190206535   0.12087003770860709   0.01428960262096088   0.1258357819093972   0.18874571653552383   0.00591102264832216   0.9087699955827645   0.4550609003324767   0.6557361540647054   0.31541201131564556   0.8801193838698916   0.41529016084485654   0.259401790704705   0.7413672207945862   0.3332247500857632   0.6666665447492519   0.666722920540872   0.9908951473552123   0.8058816452405344   0.6962458535805756   0.3946769256090145   0.014407566225027651   0.837056536972164   0.6370047237123287   0.9126806637069492   0.8935375285164205   0.8227669343512031   0.5111689418029316   0.7239349471714254   0.8876265058680984   0.9139969387684386   0.0561080414704549   0.06819879310672   0.5722144945524529   0.03387755489854696   0.6408178806255984   0.808797002402015   0.8308472737578666   0.7006528048127838   0.9741513358763464   0.14207408186114304   0.8399521264026544   0.8947711595722493   0.2779054822957709   0.7473971562521285   0.8255445601776267   0.05771462260008533   0.6409007585834421   0.8347164925451793   0.9320070316612061   0.23494768824888224   0.12973181678051052   0.11078154537375391
0.044380525793107736   0.3209507494804436   0.07362377531005564   0.04258275226703391   0.47216603124065487   0.2870731945818967   0.43280589468445724   0.23378574986501888   0.6413187574827882   0.5864203897691129   0.45865455880811085   0.09171166800387583   0.8013666310801338   0.6916492301968636   0.18074907651233993   0.3443145117517473   0.9758220709025072   0.6339346075967783   0.5398483179288978   0.509598019206568   0.043815039241301   0.39898691934789604   0.41011650114838727   0.3988164738328141   0.9994345134481932   0.07803616986745242   0.3364927258383317   0.3562337215657802   0.5272684822075384   0.7909629752855557   0.9036868311538744   0.12244797170076133   0.8859497247247502   0.20454258551644283   0.44503227234576354   0.030736303696885504   0.0845830936446163   0.5128933553195792   0.26428319583342363   0.6864217919451382   0.10876102274210915   0.8789587477228009   0.7244348779045258   0.17682377273857014   0.06494598350080814   0.4799718283749049   0.31431837675613855   0.778007298905756   0.06551147005261489   0.4019356585074525   0.9778256509178069   0.42177357733997584   0.5382429878450765   0.6109726832218967   0.0741388197639325   0.2993256056392145   0.6522932631203263   0.4064300977054539   0.629106547418169   0.268589301942329   0.5677101694757101   0.8935367423858747   0.3648233515847453   0.5821675099971908
0.4589491467336009   0.014577994663073713   0.6403884736802196   0.40534373725862066   0.3940031632327927   0.5346061662881688   0.326070096924081   0.6273364383528647   0.32849169318017785   0.13267050778071635   0.34824444600627413   0.20556286101288884   0.7902487053351014   0.5216978245588196   0.27410562624234164   0.9062372553736744   0.13795544221477501   0.11526772685336573   0.6449990788241726   0.6376479534313454   0.570245272739065   0.22173098446749107   0.28017572723942735   0.05548044343415454   0.1112961260054641   0.20715298980441735   0.6397872535592077   0.6501367061755339   0.7172929627726714   0.6725468235162485   0.3137171566351268   0.022800267822669213   0.3888012695924935   0.5398763157355322   0.9654727106288526   0.8172374068097804   0.5985525642573921   0.018178491176712597   0.6913670843865111   0.911000151436106   0.46059712204261716   0.9029107643233468   0.046368005562338346   0.2733521980047607   0.8903518493035522   0.6811797798558558   0.766192278322911   0.21787175457060615   0.779055723298088   0.47402679005143844   0.12640502476370324   0.5677350483950723   0.06176276052541669   0.8014799665351899   0.8126878681285764   0.5449347805724031   0.6729614909329231   0.2616036507996577   0.8472151574997238   0.7276973737626227   0.074408926675531   0.24342515962294511   0.15584807311321278   0.8166972223265166
0.6138118046329138   0.3405143952995982   0.10948006755087443   0.5433450243217559   0.7234599553293617   0.6593346154437424   0.3432877892279634   0.3254732697511498   0.9444042320312737   0.18530782539230398   0.21688276446426016   0.7577382213560775   0.8826414715058569   0.38382785885711407   0.40419489633568373   0.2128034407836745   0.2096799805729338   0.12222420805745636   0.55697973883596   0.4851060670210518   0.1352710538974028   0.8787990484345113   0.40113166572274717   0.6684088446945352   0.5214592492644889   0.538284653134913   0.2916515981718727   0.12506382037277922   0.7979992939351273   0.8789500376911706   0.9483638089439093   0.7995905506216294   0.8535950619038536   0.6936422122988666   0.7314810444796491   0.04185232926555184   0.9709535903979966   0.30981435344175257   0.3272861481439654   0.8290488884818773   0.7612736098250628   0.18759014538429622   0.7703064093080055   0.34394282146082555   0.62600255592766   0.30879109694978496   0.36917474358525837   0.6755339767662903   0.10454330666317106   0.770506443814872   0.07752314541338563   0.5504701563935112   0.3065440127280439   0.8915564061237014   0.12915933646947633   0.7508796057718818   0.45294895082419034   0.19791419382483472   0.3976782919898272   0.7090272765063299   0.48199536042619373   0.8880998403830821   0.07039214384586177   0.8799783880244526
0.720721750601131   0.7005096949987859   0.30008573453785625   0.536035566563627   0.09471919467347101   0.39171859804900094   0.9309109909525979   0.8605015897973367   0.9901758880103   0.621212154234129   0.8533878455392123   0.3100314334038255   0.6836318752822561   0.7296557481104277   0.724228509069736   0.5591518276319437   0.23068292445806576   0.531741554285593   0.3265502170799088   0.8501245511256137   0.748687564031872   0.6436417139025108   0.25615807323404705   0.9701461631011611   0.02796581343074103   0.9431320189037249   0.9560723386961908   0.43411059653753403   0.93324661875727   0.5514134208547239   0.025161347743592816   0.5736090067401974   0.9430707307469701   0.9302012666205949   0.1717735022043805   0.2635775733363719   0.259438855464714   0.2005455185101672   0.4475449931346445   0.7044257457044282   0.028755931006648233   0.6688039642245742   0.12099477605473574   0.8543011945788145   0.2800683669747762   0.025162250322063425   0.8648367028206887   0.8841550314776534   0.2521025535440352   0.08203023141833854   0.908764364124498   0.4500444349401193   0.31885593478676516   0.5306168105636146   0.8836030163809051   0.8764354281999219   0.3757852040397951   0.6004155439430198   0.7118295141765246   0.61285785486355   0.11634634857508108   0.39987002543285255   0.2642845210418801   0.9084321091591218
0.08759041756843285   0.7310660612082783   0.14328974498714436   0.05413091458030732   0.8075220505936567   0.7059038108862149   0.27845304216645567   0.16997588310265394   0.5554194970496215   0.6238735794678764   0.36968867804195765   0.7199314481625346   0.23656356226285627   0.09325676890426171   0.4860856616610525   0.8434960199626127   0.8607783582230611   0.49284122496124194   0.7742561474845279   0.23063816509906268   0.7444320096479801   0.09297119952838939   0.5099716264426478   0.32220605593994084   0.6568415920795473   0.36190513832011106   0.3666818814555034   0.26807514135963356   0.8493195414858906   0.6560013274338962   0.08822883928904776   0.0980992582569796   0.2939000444362692   0.03212774796601985   0.7185401612470901   0.378167810094445   0.05733648217341292   0.9388709790617581   0.2324544995860376   0.5346717901318323   0.19655812395035172   0.4460297541005162   0.4581983521015097   0.3040336250327696   0.4521261143023716   0.3530585545721268   0.948226725658862   0.9818275690928288   0.7952845222228243   0.9911534162520157   0.5815448442033585   0.7137524277331951   0.9459649807369337   0.33515208881811953   0.49331600491431077   0.6156531694762156   0.6520649363006645   0.30302434085209967   0.7747758436672206   0.23748535938177062   0.5947284541272516   0.3641533617903415   0.542321344081183   0.7028135692499383
0.3981703301768999   0.9181236076898254   0.08412299197967336   0.3987799442171687   0.9460442158745282   0.5650650531176985   0.1358962663208114   0.41695237512433997   0.1507596936517039   0.5739116368656828   0.5543514221174528   0.7031999473911448   0.2047947129147702   0.2387595480475633   0.06103541720314207   0.08754677791492921   0.5527297766141057   0.9357352071954637   0.2862595735359214   0.8500614185331586   0.9580013224868541   0.5715818454051221   0.7439382294547383   0.14724784928322027   0.5598309923099541   0.6534582377152968   0.6598152374750649   0.7484679050660515   0.6137867764354259   0.08839318459759828   0.5239189711542536   0.3315155299417116   0.46302708278372195   0.5144815477319155   0.9695675490368006   0.6283155825505667   0.25823236986895176   0.2757219996843522   0.9085321318336586   0.5407688046356376   0.7055025932548461   0.3399867924888885   0.6222725582977372   0.690707386102479   0.747501270767992   0.7684049470837664   0.8783343288429989   0.5434595368192587   0.18767027845803785   0.11494670936846958   0.21851909136793402   0.7949916317532072   0.573883502022612   0.026553524770871303   0.6946001202136804   0.4634761018114956   0.11085641923888996   0.5120719770389558   0.7250325711768798   0.8351605192609288   0.8526240493699382   0.23634997735460367   0.8165004393432213   0.2943917146252913
0.1471214561150921   0.8963631848657152   0.194227881045484   0.6036843285228123   0.3996201853471001   0.12795823778194876   0.31589355220248505   0.060224791703553625   0.21194990688906223   0.013011528413479172   0.09737446083455105   0.26523315995034646   0.6380664048664503   0.9864580036426078   0.4027743406208706   0.8017570581388508   0.5272099856275603   0.47438602660365203   0.6777417694439908   0.966596538877922   0.6745859362576221   0.23803604924904836   0.8612413301007695   0.6722048242526306   0.52746448014253   0.3416728643833332   0.6670134490552856   0.06852049572981833   0.12784429479542997   0.21371462660138446   0.3511198968528005   0.00829570402626471   0.9158943879063677   0.20070309818790527   0.25374543601824945   0.7430625440759182   0.27782798303991746   0.21424509454529742   0.8509710953973788   0.9413054859370674   0.7506179974123571   0.7398590679416454   0.1732293259533881   0.9747089470591455   0.07603206115473503   0.501823018692597   0.31198799585261855   0.3025041228065148   0.548567581012205   0.1601501543092638   0.644974546797333   0.23398362707669645   0.42072328621677507   0.9464355277078793   0.29385464994453253   0.22568792305043175   0.5048288983104073   0.7457324295199741   0.04010921392628311   0.4826253789745135   0.22700091527048985   0.5314873349746767   0.18913811852890425   0.5413198930374461
0.4763829178581327   0.7916282670330312   0.015908792575516147   0.5666109459783006   0.4003508567033977   0.28980524834043425   0.7039207967228975   0.2641068231717858   0.8517832756911927   0.12965509403117048   0.05894624992556455   0.030123196095089337   0.43105998947441765   0.18321956632329112   0.765091599981032   0.8044352730446576   0.9262310911640104   0.437487136803317   0.7249823860547489   0.3218098940701441   0.6992301758935204   0.9059998018286404   0.5358442675258447   0.780490001032698   0.22284725803538777   0.1143715347956091   0.5199354749503285   0.21387905505439742   0.8224964013319901   0.8245662864551748   0.8160146782274309   0.9497722318826116   0.9707131256407974   0.6949111924240043   0.7570684283018664   0.9196490357875223   0.5396531361663798   0.5116916261007133   0.9919768283208343   0.1152137627428647   0.6134220450023694   0.07420448929739619   0.2669944422660855   0.7934038686727206   0.914191869108849   0.1682046874687558   0.7311501747402408   0.012913867640022586   0.6913446110734612   0.0538331526731467   0.21121469978991234   0.7990348125856251   0.8688482097414711   0.22926686621797188   0.3952000215624814   0.8492625807030135   0.8981350841006738   0.5343556737939675   0.6381315932606151   0.9296135449154912   0.35848194793429394   0.022664047693254294   0.6461547649397806   0.8143997821726265
0.7450599029319245   0.9484595583958582   0.3791603226736952   0.020995913499905927   0.8308680338230755   0.7802548709271023   0.6480101479334544   0.008082045859883341   0.1395234227496143   0.7264217182539556   0.43679544814354204   0.20904723327425817   0.2706752130081432   0.4971548520359837   0.04159542658106061   0.35978465257124465   0.37254012890746946   0.9627991782420162   0.40346383332044555   0.4301711076557534   0.014058180973175504   0.9401351305487619   0.7573090683806649   0.6157713254831269   0.268998278041251   0.9916755721529038   0.37814874570696966   0.5947754119832209   0.4381302442181755   0.21142070122580148   0.7301385977735153   0.5866933661233376   0.2986068214685612   0.4849989829718459   0.29334314962997327   0.3776461328490794   0.027931608460418013   0.9878441309358622   0.25174772304891263   0.017861480277834758   0.6553914795529485   0.02504495269384597   0.8482838897284671   0.5876903726220813   0.6413332985797731   0.08490982214508407   0.09097482134780221   0.9719190471389545   0.3723350205385221   0.09323424999218027   0.7128260756408326   0.37714363515573357   0.9342047763203466   0.8818135487663787   0.9826874778673172   0.790450269032396   0.6355979548517854   0.3968145657945329   0.689344328237344   0.4128041361833166   0.6076663463913674   0.40897043485867074   0.43759660518843135   0.39494265590548183
0.9522748668384188   0.38392548216482475   0.5893127154599642   0.8072522832834005   0.3109415682586457   0.29901566001974067   0.49833789411216206   0.835333236144446   0.9386065477201236   0.20578141002756042   0.7855118184713294   0.4581896009887124   0.004401771399777123   0.32396786126118166   0.8028243406040122   0.6677393319563164   0.36880381654799177   0.9271532954666487   0.11348001236666824   0.25493519577299983   0.7611374701566244   0.518182860607978   0.6758834071782369   0.859992539867518   0.8088626033182056   0.13425737844315325   0.08657069171827263   0.052740256584117594   0.49792103505955987   0.8352417184234125   0.5882327976061106   0.21740702043967164   0.5593144873394362   0.6294603083958521   0.802720979134781   0.7592174194509592   0.5549127159396591   0.3054924471346705   0.9998966385307688   0.09147808749464281   0.1861088993916673   0.37833915166802173   0.8864166261641006   0.836542891721643   0.4249714292350429   0.8601562910600438   0.2105332189858637   0.9765503518541249   0.6161088259168374   0.7258989126168905   0.12396252726759106   0.9238100952700073   0.11818779085727746   0.8906571941934779   0.5357297296614805   0.7064030748303357   0.5588733035178413   0.2611968857976258   0.7330087505266994   0.9471856553793765   0.003960587578182224   0.9557044386629553   0.7331121119959306   0.8557075678847337
0.8178516881865149   0.5773652869949335   0.84669548583183   0.019164676163090685   0.392880258951472   0.7172089959348898   0.6361622668459663   0.04261432430896578   0.7767714330346347   0.9913100833179993   0.5121997395783753   0.11880422903895847   0.6585836421773572   0.10065288912452137   0.9764700099168948   0.4124011542086228   0.09971033865951598   0.8394560033268955   0.24346125939019536   0.46521549882924634   0.09574975108133375   0.8837515646639402   0.5103491473942647   0.6095079309445127   0.27789806289481883   0.3063862776690067   0.6636536615624348   0.590343254781422   0.8850178039433468   0.5891772817341169   0.027491394716468436   0.5477289304724562   0.10824637090871211   0.5978671984161176   0.5152916551380932   0.42892470143349776   0.4496627287313549   0.4972143092915962   0.5388216452211984   0.016523547224874972   0.34995239007183887   0.6577583059647006   0.29536038583100305   0.5513080483956286   0.25420263899050516   0.7740067413007604   0.7850112384367383   0.9418001174511159   0.9763045760956863   0.4676204636317537   0.12135757687430351   0.35145686266969395   0.09128677215233949   0.8784431818976368   0.09386618215783508   0.8037279321972377   0.9830404012436273   0.28057598348151924   0.5785745270197419   0.37480323076373995   0.5333776725122725   0.783361674189923   0.0397528817985435   0.35827968353886497
0.18342528244043363   0.12560336822522236   0.7443924959675404   0.8069716351432363   0.9292226434499286   0.351596626924462   0.9593812575308022   0.8651715176921204   0.9529180673542422   0.8839761632927082   0.8380236806564987   0.5137146550224264   0.8616312952019027   0.0055329813950714705   0.7441574984986635   0.7099867228251887   0.8785908939582753   0.7249569979135523   0.16558297147892168   0.3351834920614488   0.3452132214460028   0.9415953237236292   0.12583008968037818   0.9769038085225838   0.16178793900556915   0.8159919554984069   0.3814375937128377   0.1699321733793475   0.23256529555564065   0.46439532857394494   0.42205633618203553   0.3047606556872271   0.2796472282013985   0.5804191652812366   0.5840326555255368   0.7910460006648007   0.41801593299949574   0.5748861838861652   0.8398751570268733   0.08105927783961189   0.5394250390412204   0.8499291859726129   0.6742921855479517   0.745875785778163   0.19421181759521766   0.9083338622489837   0.5484620958675734   0.7689719772555793   0.03242387858964851   0.0923419067505768   0.16702450215473572   0.5990398038762318   0.7998585830340078   0.6279465781766319   0.7449681659727002   0.29427914818900464   0.5202113548326094   0.04752741289539521   0.1609355104471633   0.503233147524204   0.10219542183311361   0.47264122900923   0.32106035342029   0.42217386968459214
0.5627703827918932   0.6227120430366171   0.6467681678723384   0.676298083906429   0.3685585651966755   0.7143781807876334   0.09830607200476495   0.9073261066508498   0.336134686607027   0.6220362740370566   0.9312815698500292   0.308286302774618   0.5362761035730191   0.9940896958604247   0.18631340387732906   0.014007154585613352   0.01606474874040977   0.9465622829650295   0.025377893430165745   0.5107740070614093   0.9138693269072962   0.47392105395579953   0.7043175400098758   0.08860013737681721   0.351098944115403   0.8512090109191824   0.057549372137537344   0.4123020534703882   0.9825403789187275   0.136830830131549   0.9592433001327724   0.5049759468195384   0.6464056923117005   0.5147945560944924   0.027961730282743166   0.1966896440449204   0.11012958873868132   0.5207048602340677   0.8416483264054141   0.18268248945930704   0.09406483999827156   0.5741425772690382   0.8162704329752484   0.6719084823978977   0.18019551309097542   0.10022152331323862   0.11195289296537263   0.5833083450210805   0.8290965689755724   0.2490125123940562   0.05440352082783528   0.1710062915506923   0.8465561900568449   0.11218168226250719   0.09516022069506289   0.6660303447311539   0.20015049774514446   0.5973871261680148   0.06719849041231972   0.4693407006862335   0.09002090900646313   0.07668226593394711   0.2255501640069056   0.2866582112269264
0.9959560690081916   0.502539688664909   0.4092797310316572   0.6147497288290287   0.8157605559172162   0.40231816535167036   0.2973268380662846   0.03144138380794823   0.9866639869416437   0.15330565295761417   0.24292331723844932   0.8604350922572559   0.14010779688479877   0.04112397069510697   0.14776309654338643   0.19440474752610204   0.9399572991396543   0.44373684452709217   0.08056460613106671   0.7250640468398686   0.8499363901331912   0.36705457859314505   0.8550144421241611   0.4384058356129421   0.8539803211249997   0.8645148899282361   0.44573471109250384   0.8236561067839133   0.03821976520778346   0.46219672457656574   0.14840787302621924   0.7922147229759652   0.05155577826613973   0.3088910716189516   0.90548455578777   0.9317796307187092   0.911447981381341   0.2677671009238446   0.7577214592443835   0.7373748831926071   0.9714906822416867   0.8240302563967524   0.6771568531133169   0.012310836352738637   0.12155429210849546   0.4569756778036073   0.8221424109891557   0.5739050007397966   0.26757397098349583   0.5924607878753713   0.37640769989665185   0.7502488939558831   0.2293542057757124   0.13026406329880552   0.2279998268704326   0.958034170979918   0.17779842750957264   0.821372991679854   0.32251527108266265   0.026254540261208843   0.2663504461282317   0.5536058907560093   0.5647938118382791   0.2888796570686017
0.29485976388654506   0.729575634359257   0.8876369587249624   0.27656882071586303   0.1733054717780496   0.2725999565556496   0.06549454773580664   0.7026638199760665   0.9057315007945538   0.6801391686802783   0.6890868478391547   0.9524149260201833   0.6763772950188414   0.5498751053814728   0.46108702096872217   0.9943807550402652   0.4985788675092687   0.7285021137016189   0.13857174988605953   0.9681262147790565   0.23222842138103703   0.1748962229456095   0.5737779380477804   0.6792465577104547   0.9373686574944919   0.4453205885863526   0.686140979322818   0.40267773699459175   0.7640631857164424   0.17272063203070298   0.6206464315870114   0.7000139170185252   0.8583316849218886   0.49258146335042463   0.9315595837478566   0.7475989909983419   0.18195438990304721   0.9427063579689519   0.4704725627791344   0.7532182359580767   0.6833755223937785   0.21420424426733298   0.3319008128930749   0.7850920211790202   0.45114710101274147   0.039308021321723466   0.7581228748452945   0.10584546346856548   0.5137784435182495   0.5939874327353709   0.07198189552247646   0.7031677264739737   0.7497152578018071   0.42126680070466793   0.45133546393546503   0.0031538094554485136   0.8913835728799185   0.9286853373542433   0.5197758801876085   0.2555548184571066   0.7094291829768713   0.9859789793852914   0.04930331740847401   0.5023365824990299
0.02605366058309278   0.7717747351179585   0.7174025045153991   0.7172445613200097   0.5749065595703513   0.732466713796235   0.9592796296701046   0.6113990978514442   0.06112811605210184   0.1384792810608641   0.8872977341476281   0.9082313713774705   0.31141285825029474   0.7172124803561962   0.4359622702121631   0.9050775619220219   0.4200292853703762   0.7885271430019529   0.9161863900245547   0.6495227434649153   0.7106001023935049   0.8025481636166615   0.8668830726160807   0.14718616096588544   0.6845464418104121   0.030773428498703036   0.14948056810068153   0.42994159964587575   0.10963988224006084   0.29830671470246806   0.19020093843057692   0.8185425017944316   0.048511766187959   0.15982743364160393   0.30290320428294876   0.9103111304169611   0.7370989079376643   0.44261495328540773   0.8669409340707857   0.00523356849493916   0.31706962256728805   0.6540878102834549   0.9507545440462309   0.3557108250300238   0.6064695201737831   0.8515396466667934   0.08387147143015031   0.2085246640641384   0.921923078363371   0.8207662181680903   0.9343909033294687   0.7785830644182626   0.8122831961233101   0.5224595034656222   0.7441899648988919   0.9600405626238311   0.7637714299353511   0.3626320698240183   0.44128676061594313   0.04972943220687   0.026672521997686827   0.9200171165386105   0.5743458265451574   0.04449586371193084
0.7096028994303988   0.26592930625515576   0.6235912824989265   0.688785038681907   0.10313337925661566   0.41438965958836244   0.5397198110687762   0.48026037461776866   0.18121030089324472   0.5936234414202721   0.6053289077393074   0.701677310199506   0.3689271047699346   0.07116393795464986   0.8611389428404155   0.7416367475756749   0.6051556748345835   0.7085318681306315   0.4198521822244724   0.6919073153688049   0.5784831528368967   0.788514751592021   0.845506355679315   0.6474114516568741   0.8688802534064979   0.5225854453368652   0.22191507318038847   0.9586264129749671   0.7657468741498822   0.10819578574850285   0.6821952621116123   0.47836603835719843   0.5845365732566375   0.5145723443282307   0.07686635437230492   0.7766887281576924   0.21560946848670293   0.44340840637358087   0.21572741153188937   0.03505198058201748   0.6104537936521194   0.7348765382429493   0.7958752293074169   0.3431446652132126   0.03197064081522275   0.9463617866509283   0.950368873628102   0.6957332135563384   0.16309038740872486   0.42377634131406305   0.7284538004477135   0.7371068005813715   0.3973435132588426   0.31558055556556025   0.0462585383361012   0.258740762224173   0.8128069400022051   0.8010082112373295   0.9693921839637962   0.4820520340664806   0.5971974715155022   0.35759980486374865   0.7536647724319069   0.44700005348446314
0.9867436778633828   0.6227232666207994   0.9577895431244899   0.10385538827125058   0.95477303704816   0.676361479969871   0.007420669496387948   0.4081221747149121   0.7916826496394351   0.2525851386558079   0.27896686904867446   0.6710153741335407   0.39433913638059254   0.9370045830902477   0.23270833071257324   0.41227461190936765   0.5815321963783874   0.13599637185291819   0.26331614674877696   0.9302225778428871   0.9843347248628852   0.7783965669891695   0.50965137431687   0.48322252435842394   0.9975910469995025   0.1556733003683702   0.5518618311923801   0.3793671360871733   0.04281800995134253   0.47931182039849923   0.5444411616959922   0.9712449613722612   0.2511353603119074   0.2267266817426913   0.26547429264731776   0.30022958723872056   0.8567962239313149   0.28972209865244364   0.03276596193474449   0.8879549753293529   0.27526402755292745   0.15372572679952545   0.7694498151859676   0.9577323974864658   0.2909293026900422   0.3753291598103559   0.2597984408690975   0.4745098731280419   0.2933382556905397   0.2196558594419857   0.7079366096767173   0.09514273704086855   0.2505202457391972   0.7403440390434864   0.16349544798072518   0.12389777566860731   0.9993848854272898   0.5136173573007952   0.8980211553334074   0.8236681884298868   0.14258866149597488   0.22389525864835155   0.865255193398663   0.9357132131005339
0.8673246339430474   0.07016953184882613   0.09580537821269541   0.977980815614068   0.5763953312530052   0.6948403720384703   0.8360069373435979   0.5034709424860262   0.2830570755624655   0.47518451259648453   0.1280703276668806   0.40832820544515763   0.03253682982326838   0.7348404735529981   0.9645748796861554   0.2844304297765503   0.03315194439597862   0.22122311625220287   0.06655372435274795   0.46076224134666355   0.8905632829000037   0.9973278576038513   0.201298530954085   0.5250490282461296   0.02323864895695632   0.9271583257550252   0.1054931527413896   0.5470682126320616   0.4468433177039511   0.23231795371655495   0.26948621539779166   0.04359727014603542   0.16378624214148557   0.7571334411200704   0.14141588773091107   0.6352690647008779   0.13124941231821718   0.022292967567072403   0.1768410080447557   0.35083863492432754   0.09809746792223857   0.8010698513148695   0.11028728369200774   0.890076393577664   0.20753418502223483   0.8037419937110183   0.9089887527379228   0.36502736533153435   0.18429553606527851   0.8765836679559931   0.8034955999965332   0.8179591526994727   0.7374522183613275   0.6442657142394381   0.5340093845987415   0.7743618825534373   0.5736659762198418   0.8871322731193677   0.3925934968678304   0.1390928178525595   0.44241656390162465   0.8648393055522953   0.2157524888230747   0.788254182928232
0.3443190959793861   0.06376945423742572   0.10546520513106698   0.898177789350568   0.13678491095715123   0.26002746052640746   0.19647645239314424   0.5331504240190337   0.9524893748918727   0.3834437925704144   0.3929808523966111   0.715191271319561   0.2150371565305453   0.7391780783309763   0.8589714677978696   0.9408293887661237   0.6413711803107035   0.8520458052116087   0.46637797093003924   0.8017365709135641   0.19895461640907883   0.9872064996593134   0.2506254821069645   0.01348238798533212   0.8546355204296927   0.9234370454218876   0.14516027697589753   0.11530459863476411   0.7178506094725415   0.6634095848954802   0.9486838245827532   0.5821541746157304   0.7653612345806687   0.2799657923250658   0.5557029721861422   0.8669629032961695   0.5503240780501235   0.5407877139940894   0.6967315043882726   0.9261335145300459   0.90895289773942   0.6887419087824809   0.23035353345823334   0.12439694361648176   0.7099982813303412   0.7015354091231675   0.9797280513512688   0.11091455563114964   0.8553627609006483   0.7780983637012798   0.8345677743753713   0.9956099569963855   0.13751215142810685   0.11468877880579963   0.8858839497926181   0.4134557823806551   0.37215091684743806   0.8347229864807338   0.33018097760647586   0.5464928790844856   0.8218268387973147   0.29393527248664436   0.6334494732182033   0.6203593645544397
0.9128739410578947   0.6051933637041635   0.40309593975996993   0.495962420937958   0.20287565972755348   0.9036579545809961   0.4233678884087011   0.38504786530680835   0.3475128988269051   0.12555959087971624   0.5888001140333298   0.3894379083104228   0.21000074739879823   0.010870812073916625   0.7029161642407118   0.9759821259297677   0.8378498305513602   0.17614782559318276   0.3727351866342359   0.4294892468452821   0.01602299175404554   0.8822125531065383   0.7392857134160327   0.8091298822908424   0.1031490506961509   0.27701918940237485   0.3361897736560627   0.31316746135288437   0.9002733909685975   0.3733612348213788   0.9128218852473616   0.9281195960460761   0.5527604921416923   0.2478016439416625   0.3240217712140318   0.5386816877356532   0.3427597447428941   0.2369308318677459   0.6211056069733201   0.5626995618058855   0.504909914191534   0.06078300627456313   0.24837042033908419   0.13321031496060343   0.48888692243748844   0.17857045316802475   0.5090847069230516   0.3240804326697611   0.3857378717413375   0.9015512637656499   0.1728949332669889   0.010912971316876722   0.48546448077274007   0.5281900289442711   0.26007304801962733   0.08279337527080069   0.9327039886310478   0.2803883850026086   0.9360512768055955   0.5441116875351475   0.5899442438881536   0.04345755313486267   0.3149456698322754   0.981412125729262
0.08503432969661966   0.9826745468602995   0.06657524949319123   0.8482018107686585   0.5961474072591313   0.8041040936922748   0.5574905425701396   0.5241213780988975   0.21040953551779373   0.9025528299266249   0.38459560930315073   0.5132084067820207   0.7249450547450537   0.3743628009823538   0.12452256128352343   0.43041503151122   0.7922410661140059   0.09397441597974523   0.18847128447792794   0.8863033439760726   0.20229682222585232   0.05051686284488256   0.8735256146456525   0.9048912182468106   0.11726249252923265   0.06784231598458303   0.8069503651524613   0.056689407478152064   0.5211150852701014   0.2637382222923082   0.24945982258232166   0.5325680293792546   0.3107055497523077   0.3611853923656833   0.864864213279171   0.019359622597233905   0.585760495007254   0.9868225913833295   0.7403416519956475   0.5889445910860139   0.7935194288932481   0.8928481754035843   0.5518703675177196   0.7026412471099414   0.5912226066673958   0.8423313125587018   0.678344752872067   0.7977500288631307   0.4739601141381631   0.7744889965741186   0.8713943877196056   0.7410606213849786   0.9528450288680617   0.5107507742818105   0.6219345651372841   0.20849259200572406   0.642139479115754   0.14956538191612714   0.7570703518581131   0.18913296940849014   0.0563789841085   0.16274279053279767   0.016728699862465675   0.6001883783224763
0.26285955521525195   0.2698946151292134   0.46485833234474616   0.8975471312125349   0.6716369485478562   0.42756330257051167   0.7865135794726792   0.09979710234940418   0.19767683440969308   0.653074305996393   0.9151191917530734   0.3587364809644255   0.2448318055416314   0.14232353171458256   0.2931846266157894   0.15024388895870144   0.6026923264258773   0.9927581497984554   0.5361142747576763   0.9611109195502113   0.5463133423173774   0.8300153592656577   0.5193855748952105   0.36092254122773504   0.28345378710212543   0.5601207441364443   0.054527242550464435   0.4633754100152001   0.6118168385542693   0.13255744156593266   0.2680136630777853   0.3635783076657959   0.4141400041445762   0.47948313556953964   0.35289447132471186   0.004841826701370412   0.16930819860294483   0.3371596038549571   0.05970984470892244   0.854597937742669   0.5666158721770674   0.3444014540565017   0.5235955699512462   0.8934870181924577   0.020302529859690048   0.514386094790844   0.004209995056035597   0.5325644769647226   0.7368487427575646   0.9542653506543995   0.9496827525055712   0.06918906694952251   0.12503190420329532   0.8217079090884669   0.6816690894277859   0.7056107592837266   0.710891900058719   0.34222477351892727   0.328774618103074   0.7007689325823562   0.5415837014557743   0.005065169663970205   0.2690647733941516   0.8461709948396873
0.9749678292787068   0.6606637156074685   0.7454692034429055   0.9526839766472296   0.9546652994190168   0.14627762081662463   0.7412592083868699   0.42011949968250695   0.21781655666145222   0.19201227016222505   0.7915764558812987   0.35093043273298447   0.09278465245815691   0.37030436107375814   0.10990736645351279   0.6453196734492579   0.3818927523994378   0.028079587554830872   0.7811327483504388   0.9445507408669017   0.8403090509436635   0.023014417890860665   0.5120679749562872   0.09837974602721446   0.8653412216649566   0.3623507022833921   0.7665987715133817   0.14569576937998488   0.9106759222459399   0.2160730814667675   0.025339563126511904   0.7255762696974779   0.6928593655844877   0.024060811304542445   0.23376310724521324   0.3746458369644935   0.6000747131263308   0.6537564502307843   0.12385574079170046   0.7293261635152356   0.21818196072689292   0.6256768626759535   0.3427229924412617   0.784775422648334   0.3778729097832294   0.6026624447850928   0.8306550174849746   0.6863956766211196   0.5125316881182728   0.24031174250170062   0.06405624597159283   0.5406999072411346   0.6018557658723329   0.024238661034933127   0.03871668284508093   0.8151236375436567   0.9089964002878452   0.0001778497303906825   0.8049535755998677   0.4404778005791632   0.3089216871615146   0.3464213994996064   0.6810978348081672   0.7111516370639276
0.09073972643462162   0.7207445368236529   0.3383748423669055   0.9263762144155936   0.7128668166513922   0.1180820920385602   0.5077198248819309   0.23998053779447404   0.20033512853311947   0.8777703495368596   0.44366357891033814   0.6992806305533394   0.5984793626607865   0.8535316885019264   0.4049468960652572   0.8841569930096826   0.6894829623729413   0.8533538387715357   0.5999933204653896   0.4436791924305195   0.3805612752114267   0.5069324392719293   0.9188954856572222   0.732527555366592   0.28982154877680505   0.7861879024482764   0.5805206432903167   0.8061513409509984   0.5769547321254128   0.6681058104097162   0.07280081840838581   0.5661708031565243   0.3766196035922934   0.7903354608728567   0.6291372394980477   0.8668901726031849   0.7781402409315069   0.9368037723709303   0.2241903434327905   0.9827331795935023   0.08865727855856562   0.08344993359939445   0.624197022967401   0.5390539871629827   0.708096003347139   0.5765174943274651   0.7053015373101787   0.8065264317963908   0.41827445457033385   0.7903295918791887   0.12478089401986195   0.0003750908453924338   0.8413197224449209   0.12222378146947246   0.05198007561147615   0.4342042876888681   0.4647001188526276   0.3318883205966158   0.42284283611342843   0.5673141150856832   0.6865598779211207   0.3950845482256856   0.19865249268063795   0.5845809354921809
0.5979025993625551   0.31163461462629116   0.5744554697132369   0.045526948329198236   0.8898065960154162   0.735117120298826   0.8691539324030583   0.23900051653280743   0.4715321414450823   0.9447875284196374   0.7443730383831962   0.23862542568741502   0.6302124190001613   0.8225637469501649   0.6923929627717201   0.8044211379985469   0.1655123001475338   0.4906754263535491   0.2695501266582917   0.2371070229128637   0.4789524222264131   0.09559087812786349   0.07089763397765372   0.6525260874206827   0.881049822863858   0.7839562635015723   0.4964421642644168   0.6069991390914845   0.9912432268484418   0.04883914320274628   0.6272882318613585   0.36799862255867705   0.5197110854033595   0.1040516147831089   0.8829151934781623   0.12937319687126206   0.8894986664031981   0.281487867832944   0.1905222307064421   0.32495205887271517   0.7239863662556644   0.7908124414793949   0.9209721040481504   0.08784503595985146   0.24503394402925122   0.6952215633515314   0.8500744700704966   0.43531894853916875   0.3639841211653932   0.9112652998499591   0.3536323058060799   0.8283198094476842   0.37274089431695134   0.8624261566472128   0.7263440739447214   0.4603211868890072   0.8530298089135919   0.7583745418641039   0.8434288804665592   0.33094799001774516   0.9635311425103937   0.4768866740311599   0.652906649760117   0.005995931145029977
0.23954477625472942   0.686074232551765   0.7319345457119667   0.9181508951851786   0.9945108322254782   0.9908526692002336   0.88186007564147   0.48283194664600976   0.630526711060085   0.07958736935027455   0.5282277698353901   0.6545121371983256   0.2577858167431336   0.21716121270306177   0.8018836958906687   0.19419095030931835   0.40475600782954174   0.4587866708389579   0.9584548154241095   0.8632429602915732   0.441224865319148   0.9818999968077979   0.3055481656639924   0.8572470291465433   0.2016800890644186   0.29582576425603296   0.5736136199520258   0.9390961339613647   0.2071692568389404   0.30497309505579934   0.6917535443105558   0.45626418731535495   0.5766425457788554   0.22538572570552481   0.16352577447516575   0.8017520501170294   0.3188567290357218   0.008224513002463038   0.3616420785844971   0.6075610998077111   0.9141007212061801   0.5494378421635051   0.4031872631603876   0.7443181395161379   0.4728758558870321   0.5675378453557072   0.09763909749639518   0.8870711103695946   0.27119576682261354   0.2717120810996742   0.5240254775443695   0.9479749764082299   0.06402650998367311   0.9667389860438749   0.8322719332338137   0.49171078909287497   0.48738396420481767   0.74135326033835   0.6687461587586478   0.6899587389758456   0.16852723516909585   0.733128747335887   0.3071040801741508   0.08239763916813451
0.2544265139629157   0.18369090517238185   0.9039168170137631   0.33807949965199663   0.7815506580758836   0.6161530598166747   0.806277719517368   0.451008389282402   0.51035489125327   0.34444097871700047   0.2822522419729986   0.5030334128741721   0.446328381269597   0.37770199267312565   0.44998030873918493   0.011322623781297114   0.9589444170647793   0.6363487323347756   0.7812341499805371   0.3213638848054515   0.7904171818956834   0.9032199849988886   0.4741300698063863   0.23896624563731703   0.5359906679327677   0.7195290798265067   0.570213252792623   0.9008867459853204   0.7544400098568841   0.10337602000983208   0.7639355332752551   0.44987835670291837   0.244085118603614   0.7589350412928316   0.48168329130225646   0.9468449438287463   0.797756737334017   0.38123304861970597   0.03170298256307153   0.9355223200474492   0.8388123202692377   0.7448843162849303   0.2504688325825345   0.6141584352419976   0.04839513837355424   0.8416643312860418   0.7763387627761482   0.3751921896046806   0.5124044704407865   0.12213525145953501   0.20612550998352513   0.4743054436193602   0.7579644605839024   0.01875923144970293   0.4421899767082701   0.024427086916441874   0.5138793419802884   0.2598241901568713   0.9605066854060136   0.07758214308769563   0.7161226046462713   0.8785911415371653   0.9288037028429421   0.1420598230402465
0.8773102843770336   0.13370682525223498   0.6783348702604076   0.5279013877982489   0.8289151460034794   0.29204249396619325   0.9019961074842594   0.15270919819356832   0.3165106755626929   0.1699072425066582   0.6958705975007342   0.6784037545742081   0.5585462149787905   0.15114801105695527   0.2536806207924642   0.6539766676577662   0.04466687299850211   0.891323820900084   0.29317393538645053   0.5763945245700706   0.3285442683522308   0.012732679362918596   0.3643702325435085   0.4343347015298241   0.4512339839751971   0.8790258541106836   0.6860353622831009   0.9064333137315752   0.6223188379717177   0.5869833601444904   0.7840392547988415   0.7537241155380069   0.3058081624090248   0.41707611763783214   0.08816865729810724   0.07532036096379877   0.7472619474302343   0.2659281065808769   0.8344880365056431   0.42134369330603255   0.7025950744317322   0.37460428568079296   0.5413141011191925   0.8449491687359619   0.3740508060795014   0.36187160631787435   0.17694386857568403   0.4106144672061378   0.9228168221043044   0.4828457522071907   0.49090850629258315   0.5041811534745626   0.3004979841325866   0.8958623920627004   0.7068692514937417   0.7504570379365557   0.9946898217235618   0.47878627442486815   0.6187005941956344   0.6751366769727569   0.24742787429332752   0.21285816784399128   0.7842125576899913   0.2537929836667244
0.5448327998615953   0.8382538821631984   0.24289845657079884   0.4088438149307625   0.17078199378209388   0.476382275845324   0.0659545879951148   0.9982293477246247   0.24796517167778953   0.9935365236381333   0.5750460817025317   0.4940481942500621   0.9474671875452029   0.09767413157543293   0.86817683020879   0.7435911563135064   0.9527773658216411   0.6188878571505647   0.24947623601315552   0.06845447934074937   0.7053494915283136   0.40602968930657346   0.4652636783231642   0.8146614956740249   0.16051669166671825   0.5677758071433752   0.2223652217523653   0.4058176807432624   0.9897346978846244   0.09139353129805111   0.1564106337572505   0.4075883330186377   0.7417695262068349   0.09785700765991782   0.5813645520547188   0.9135401387685756   0.7943023386616319   0.00018287608448488155   0.7131877218459289   0.1699489824550693   0.8415249728399908   0.3812950189339201   0.4637114858327734   0.10149450311431991   0.1361754813116773   0.9752653296273467   0.9984478075096093   0.286833007440295   0.975658789644959   0.4074895224839715   0.776082585757244   0.8810153266970325   0.9859240917603347   0.3160959911859204   0.6196719519999934   0.47342699367839486   0.2441545655534998   0.21823898352600257   0.038307399945274545   0.5598868549098193   0.4498522268918678   0.21805610744151768   0.3251196780993456   0.38993787245475
0.6083272540518769   0.8367610885075976   0.8614081922665723   0.28844336934043   0.47215177274019965   0.861495758880251   0.862960384756963   0.001610361900135064   0.49649298309524065   0.45400623639627946   0.08687779899971908   0.1205950352031025   0.510568891334906   0.13791024521035905   0.46720584699972567   0.6471680415247076   0.26641432578140617   0.9196712616843564   0.4288984470544511   0.0872811866148884   0.8165620988895383   0.7016151542428388   0.10377876895510547   0.6973433141601384   0.20823484483766136   0.8648540657352412   0.24237057668853323   0.4088999448197084   0.7360830720974617   0.003358306854990253   0.3794101919315702   0.40728958291957335   0.23959008900222106   0.5493520704587108   0.2925323929318512   0.28669454771647085   0.7290211976673151   0.41144182524835177   0.8253265459321255   0.6395265061917632   0.46260687188590893   0.49177056356399534   0.3964280988776744   0.5522453195768748   0.6460447729963706   0.7901554093211566   0.2926493299225689   0.8549020054167363   0.4378099281587092   0.9253013435859153   0.050278753234035696   0.44600206059702796   0.7017268560612476   0.9219430367309251   0.6708685613024654   0.038712477677454615   0.4621367670590265   0.3725909662722143   0.3783361683706143   0.7520179299609838   0.7331155693917114   0.9611491410238625   0.5530096224384888   0.11249142376922056
0.27050869750580253   0.46937857745986716   0.1565815235608144   0.5602461041923458   0.6244639245094319   0.6792231681387106   0.8639321936382455   0.7053440987756094   0.18665399635072266   0.7539218245527953   0.8136534404042097   0.2593420381785814   0.4849271402894751   0.8319787878218702   0.1427848791017443   0.2206295605011268   0.02279037323044857   0.4593878215496559   0.76444871073113   0.46861163054014304   0.2896748038387371   0.4982386805257934   0.21143908829264121   0.3561202067709225   0.019166106332934613   0.028860103065926235   0.054857564731826826   0.7958741025785767   0.3947021818235027   0.3496369349272156   0.19092537109358135   0.09053000380296736   0.20804818547278003   0.5957151103744203   0.3772719306893716   0.8311879656243859   0.7231210451833049   0.7637363225525501   0.23448705158762725   0.6105584051232591   0.7003306719528564   0.30434850100289423   0.47003834085649726   0.14194677458311605   0.41065586811411925   0.8061098204771008   0.258599252563856   0.7858265678121935   0.3914897617811846   0.7772497174111745   0.2037416878320292   0.9899524652336168   0.996787579957682   0.42761278248395895   0.012816316738447847   0.8994224614306494   0.7887393944849019   0.8318976721095387   0.6355443860490763   0.06823449580626352   0.06561834930159698   0.06816134955698853   0.401057334461449   0.4576760906830044
0.3652876773487406   0.7638128485540944   0.9310189936049518   0.31572931609988836   0.9546318092346214   0.9577030280769935   0.6724197410410957   0.5299027482876948   0.5631420474534368   0.18045331066581896   0.4686780532090665   0.539950283054078   0.5663544674957548   0.75284052818186   0.4558617364706187   0.6405278216234286   0.777615073010853   0.9209428560723213   0.8203173504215424   0.5722933258171651   0.7119967237092559   0.8527815065153328   0.4192600159600934   0.11461723513416062   0.34670904636051536   0.08896865796123848   0.48824102235514166   0.7988879190342723   0.392077237125894   0.13126562988424498   0.815821281314046   0.26898517074657746   0.8289351896724572   0.950812319218426   0.3471432281049794   0.7290348876924995   0.26258072217670236   0.19797179103656604   0.8912814916343608   0.0885070660690709   0.48496564916584944   0.2770289349642447   0.07096414121281833   0.5162137402519058   0.7729689254565935   0.4242474284489119   0.6517041252527249   0.40159650511774525   0.4262598790960781   0.3352787704876734   0.16346310289758328   0.602708586083473   0.0341826419701841   0.20401314060342843   0.34764182158353735   0.33372341533689553   0.2052474522977269   0.2532008213850024   0.0004985934785579455   0.6046885276443961   0.9426667301210245   0.05522903034843637   0.10921710184419721   0.5161814615753252
0.4577010809551751   0.7782000953841917   0.03825296063137888   0.9999677213234193   0.6847321554985817   0.35395266693527977   0.386548835378654   0.598371216205674   0.2584722764025036   0.018673896447606385   0.22308573248107066   0.9956626301222011   0.22428963443231947   0.814660755844178   0.8754439108975334   0.6619392147853056   0.019042182134592595   0.5614599344591755   0.8749453174189754   0.05725068714090954   0.07637545201356807   0.5062309041107392   0.7657282155747782   0.5410692255655843   0.618674371058393   0.7280308087265475   0.7274752549433993   0.5411015042421651   0.9339422155598113   0.37407814179126775   0.34092641956474534   0.9427302880364911   0.6754699391573077   0.35540424534366133   0.11784068708367466   0.9470676579142899   0.4511803047249882   0.5407434894994834   0.24239677618614133   0.28512844312898433   0.43213812259039563   0.9792835550403078   0.36745145876716595   0.22787775598807478   0.3557626705768276   0.47305265092956866   0.6017232431923878   0.6868085304224903   0.7370882995184346   0.7450218422030211   0.8742479882489885   0.1457070261803253   0.8031460839586233   0.3709437004117534   0.5333215686842432   0.2029767381438343   0.12767614480131556   0.015539455068092064   0.4154808816005685   0.25590908022954434   0.6764958400763273   0.4747959655686087   0.17308410541442718   0.9707806371005601
0.24435771748593169   0.49551241052830086   0.8056326466472612   0.7429028811124853   0.8885950469091041   0.022459759598732226   0.2039094034548734   0.05609435068999484   0.15150674739066952   0.2774379173957111   0.3296614152058849   0.9103873245096695   0.3483606634320462   0.9064942169839577   0.7963398465216417   0.7074105863658352   0.22068451863073066   0.8909547619158656   0.3808589649210732   0.45150150613629086   0.5441886785544033   0.41615879634725694   0.207774859506646   0.48072086903573086   0.2998309610684716   0.9206463858189561   0.4021422128593848   0.7378179879232456   0.4112359141593675   0.8981866262202238   0.19823280940451138   0.6817236372332508   0.259729166768698   0.6207487088245127   0.8685713941986265   0.7713363127235813   0.9113685033366518   0.7142544918405551   0.07223154767698475   0.063925726357746   0.6906839847059212   0.8232997299246895   0.6913725827559116   0.6124242202214552   0.14649530615151782   0.4071409335774325   0.4835977232492656   0.13170335118572427   0.8466643450830462   0.4864945477584764   0.08145551038988079   0.3938853632624787   0.43542843092367867   0.5883079215382525   0.8832227009853694   0.7121617260292279   0.1756992641549807   0.9675592127137398   0.014651306786742951   0.9408254133056466   0.2643307608183289   0.25330472087318473   0.9424197591097582   0.8768996869479007
0.5736467761124078   0.4300049909484953   0.2510471763538466   0.2644754667264455   0.42715146996089   0.022864057371062806   0.767449453104581   0.13277211554072124   0.5804871248778438   0.5363695096125864   0.6859939427147003   0.7388867522782426   0.1450586939541651   0.9480615880743338   0.8027712417293309   0.026725026249014686   0.9693594297991844   0.9805023753605941   0.7881199349425879   0.08589961294336804   0.7050286689808555   0.7271976544874094   0.8457001758328297   0.20899992599546738   0.1313818928684477   0.2971926635389141   0.5946529994789831   0.9445244592690218   0.7042304229075578   0.27432860616785126   0.8272035463744021   0.8117523437283006   0.12374329802971396   0.7379590965552649   0.14120960365970175   0.07286559145005801   0.9786846040755489   0.789897508480931   0.3384383619303709   0.04614056520104333   0.009325174276364472   0.809395133120337   0.550318426987783   0.9602409522576753   0.304296505295509   0.08219747863292752   0.7046182511549534   0.7512410262622079   0.1729146124270613   0.7850048150940134   0.10996525167597022   0.8067165669931861   0.4686841895195036   0.5106762089261622   0.2827617053015682   0.9949642232648854   0.3449408914897896   0.7727171123708972   0.14155210164186646   0.9220986318148274   0.36625628741424077   0.9828196038899663   0.8031137397114956   0.8759580666137841
0.3569311131378763   0.17342447076962936   0.25279531272371253   0.9157171143561088   0.052634607842367294   0.09122699213670182   0.5481770615687592   0.16447608809390088   0.879719995415306   0.3062221770426884   0.438211809892789   0.35775952110071485   0.4110358058958024   0.7955459681165262   0.15545010459122077   0.36279529783582937   0.06609491440601278   0.022828855745628984   0.013898002949354336   0.44069666602100194   0.699838626991772   0.040009251855662724   0.2107842632378588   0.5647385994072178   0.34290751385389573   0.8665847810860333   0.9579889505141462   0.649021485051109   0.29027290601152844   0.7753577889493315   0.40981188894538706   0.4845453969572081   0.41055291059622245   0.46913561190664316   0.971600079052598   0.12678587585649329   0.9995171047004201   0.6735896437901169   0.8161499744613773   0.763990578020664   0.9334221902944072   0.6507607880444879   0.802251971512023   0.323293911999662   0.23358356330263524   0.6107515361888252   0.5914677082741642   0.7585553125924441   0.8906760494487395   0.7441667551027918   0.6334787577600178   0.10953382754133519   0.600403143437211   0.9688089661534602   0.22366686881463083   0.6249884305841271   0.18985023284098856   0.49967335424681714   0.2520667897620328   0.4982025547276338   0.19033312814056852   0.8260837104567003   0.4359168153006555   0.7342119767069699
0.25691093784616126   0.17532292241221234   0.6336648437886325   0.4109180647073079   0.023327374543526038   0.5645713862233872   0.04219713551446842   0.6523627521148637   0.13265132509478655   0.8204046311205954   0.4087183777544506   0.5428289245735285   0.5322481816575755   0.851595664967135   0.18505150893981973   0.9178404939894015   0.3423979488165869   0.35192231072031793   0.9329847191777869   0.4196379392617676   0.1520648206760184   0.5258386002636177   0.49706790387713146   0.6854259625547977   0.8951538828298572   0.3505156778514053   0.8634030600884989   0.2745078978474898   0.8718265082863311   0.7859442916280182   0.8212059245740305   0.6221451457326261   0.7391751831915445   0.9655396605074228   0.41248754681957994   0.07931622115909756   0.20692700153396903   0.11394399554028775   0.2274360378797602   0.16147572716969613   0.8645290527173821   0.7620216848199698   0.2944513187019732   0.7418377879079285   0.7124642320413637   0.23618308455635215   0.7973834148248418   0.056411825353130766   0.8173103492115066   0.8856674067049468   0.9339803547363429   0.781903927505641   0.9454838409251755   0.09972311507692866   0.11277443016231241   0.15975878177301486   0.20630865773363088   0.13418345456950584   0.7002868833427325   0.0804425606139173   0.9993816561996619   0.02023945902921808   0.4728508454629723   0.9189668334442211
0.13485260348227976   0.25821777420924824   0.17839952676099907   0.1771290455362927   0.42238837144091607   0.022034689652896088   0.3810161119361573   0.12071722018316192   0.6050780222294095   0.13636728294794925   0.4470357571998144   0.33881329267752097   0.6595941813042341   0.0366441678710206   0.334261327037502   0.1790545109045061   0.45328552357060314   0.9024607133015148   0.6339744436947695   0.09861195029058882   0.4539038673709413   0.8822212542722967   0.16112359823179723   0.17964511684636764   0.31905126388866156   0.6240034800630484   0.9827240714707981   0.00251607131007495   0.8966628924477454   0.6019687904101524   0.6017079595346408   0.881798851126913   0.291584870218336   0.4656015074622031   0.15467220233482643   0.542985558449392   0.6319906889141019   0.4289573395911825   0.8204108752973244   0.3639310475448859   0.17870516534349878   0.5264966262896678   0.18643643160255488   0.26531909725429714   0.7248012979725574   0.6442753720173711   0.025312833370757643   0.08567398040792949   0.4057500340838959   0.020271891954322607   0.04258876189995949   0.08315790909785453   0.5090871416361504   0.4183031015441703   0.4408808023653186   0.2013590579709415   0.21750227141781445   0.9527015940819672   0.2862086000304922   0.6583734995215494   0.5855115825037125   0.5237442544907847   0.46579772473316783   0.2944424519766635
0.40680641716021376   0.997247628201117   0.279361293130613   0.029123354722366386   0.6820051191876563   0.35297225618374595   0.2540484597598553   0.9434493743144369   0.27625508510376034   0.33270036422942334   0.21145969785989582   0.8602914652165824   0.7671679434676099   0.914397262685253   0.7705788954945771   0.6589324072456408   0.5496656720497954   0.9616956686032859   0.48437029546408494   0.0005589077240913949   0.964154089546083   0.43795141411250116   0.01857257073091713   0.7061164557474279   0.5573476723858692   0.4407037859113842   0.7392112776003041   0.6769931010250615   0.875342553198213   0.08773152972763827   0.48516281784044885   0.7335437267106246   0.5990874680944526   0.7550311654982149   0.2737031199805531   0.8732522614940422   0.8319195246268427   0.8406339028129619   0.5031242244859758   0.2143198542484014   0.2822538525770472   0.878938234209676   0.018753929021890926   0.21376094652431   0.3180997630309643   0.4409868200971748   0.00018135829097379514   0.5076444907768821   0.7607520906450951   0.0002830341857906105   0.2609700806906696   0.8306513897518206   0.8854095374468822   0.9125515044581524   0.7758072628502207   0.09710766304119602   0.2863220693524296   0.1575203389599374   0.5021041428696676   0.22385540154715378   0.45440254472558694   0.3168864361469755   0.9989799183836918   0.00953554729875238
0.1721486921485397   0.4379482019372995   0.9802259893618009   0.7957746007744424   0.8540489291175754   0.9969613818401247   0.9800446310708271   0.2881301099975603   0.09329683847248027   0.996678347654334   0.7190745503801574   0.45747872024573966   0.20788730102559808   0.08412684319618173   0.9432672875299367   0.36037105720454365   0.9215652316731685   0.9266065042362444   0.441163144660269   0.13651565565738985   0.46716268694758156   0.6097200680892688   0.4421832262765772   0.1269801083586375   0.2950139947990419   0.17177186615196935   0.4619572369147763   0.3312055075841951   0.4409650656814665   0.17481048431184468   0.4819126058439492   0.04307539758663483   0.3476682272089862   0.1781321366575106   0.7628380554637917   0.5855966773408952   0.1397809261833881   0.09400529346132888   0.819570767933855   0.22522562013635153   0.21821569451021963   0.16739878922508453   0.37840762327358596   0.08870996447896168   0.751053007562638   0.5576787211358157   0.9362243969970088   0.9617298561203242   0.4560390127635962   0.38590685498384636   0.4742671600822324   0.630524348536129   0.015073947082129738   0.21109637067200168   0.9923545542382832   0.5874489509494942   0.6674057198731436   0.03296423401449106   0.2295164987744915   0.0018522736085990863   0.5276247936897555   0.9389589405531622   0.4099457308406365   0.7766266534722476
0.3094090991795358   0.7715601513280776   0.03153810756705056   0.6879166889932858   0.5583560916168977   0.21388143019226197   0.09531371057004183   0.7261868328729617   0.1023170788533015   0.8279745752084157   0.6210465504878094   0.09566248433683258   0.08724313177117177   0.616878204536414   0.6286919962495262   0.5082135333873383   0.41983741189802826   0.5839139705219228   0.39917549747503467   0.5063612597787392   0.8922126182082728   0.6449550299687606   0.9892297666343981   0.7297346063064917   0.582803519028737   0.873394878640683   0.9576916590673475   0.04181791731320581   0.024447427411839282   0.6595134484484211   0.8623779484973058   0.3156310844402441   0.9221303485585378   0.8315388732400054   0.24133139800949638   0.21996860010341157   0.834887216787366   0.21466066870359152   0.6126394017599702   0.7117550667160732   0.4150498048893378   0.6307466981816686   0.21346390428493553   0.20539380693733403   0.5228371866810649   0.985791668212908   0.22423413765053737   0.4756592006308423   0.940033667652328   0.11239678957222492   0.2665424785831898   0.43384128331763655   0.9155862402404887   0.45288334112380385   0.40416453008588404   0.1182101988773924   0.9934558916819509   0.6213444678837984   0.16283313207638767   0.8982415987739808   0.1585686748945849   0.40668379918020686   0.5501937303164175   0.18648653205790758
0.7435188700052471   0.7759371009985382   0.33672982603148194   0.9810927251205735   0.22068168332418214   0.7901454327856302   0.11249568838094455   0.5054335244897312   0.28064801567185416   0.6777486432134053   0.8459532097977548   0.07159224117209466   0.3650617754313655   0.22486530208960145   0.4417886797118707   0.9533820422947022   0.37160588374941456   0.603520834205803   0.278955547635483   0.05514044352072143   0.21303720885482966   0.19683703502559627   0.7287618173190655   0.8686539114628139   0.46951833884958255   0.42089993402705805   0.39203199128758365   0.8875611863422403   0.24883665552540038   0.6307545012414278   0.2795363029066391   0.3821276618525091   0.9681886398535462   0.9530058580280225   0.4335830931088844   0.31053542068041445   0.6031268644221807   0.7281405559384211   0.9917944133970137   0.3571533783857122   0.23152098067276614   0.12461972173261797   0.7128388657615307   0.30201293486499076   0.01848377181793646   0.9277826867070217   0.984077048442465   0.4333590234021769   0.5489654329683539   0.5068827526799636   0.5920450571548814   0.5457978370599366   0.3001287774429535   0.8761282514385358   0.3125087542482423   0.1636701752074275   0.3319401375894073   0.9231223934105133   0.878925661139358   0.853134754527013   0.7288132731672267   0.1949818374720922   0.8871312477423443   0.49598137614130083
0.4972922924944605   0.07036211573947421   0.17429238198081368   0.19396844127631008   0.4788085206765241   0.1425794290324525   0.19021533353834866   0.7606094178741332   0.9298430877081701   0.6356966763524888   0.5981702763834673   0.21481158081419657   0.6297143102652166   0.759568424913953   0.28566152213522494   0.05114140560676908   0.29777417267580925   0.8364460315034398   0.406735860995867   0.19800665107975604   0.5689608995085826   0.6414641940313476   0.5196046132535227   0.7020252749384552   0.07166860701412209   0.5711020782918734   0.34531223127270905   0.5080568336621452   0.592860086337598   0.4285226492594209   0.1550968977343604   0.747447415788012   0.6630169986294279   0.792825972906932   0.5569266213508931   0.5326358349738154   0.03330268836421133   0.033257547992979   0.27126509921566816   0.48149442936704634   0.735528515688402   0.1968115164895392   0.8645292382198011   0.28348777828729027   0.1665676161798195   0.5553473224581916   0.3449246249662784   0.5814625033488351   0.09489900916569742   0.9842452441663182   0.9996123936935694   0.07340566968668992   0.5020389228280994   0.5557225949068972   0.8445154959592089   0.32595825389867794   0.8390219241986715   0.7628966219999652   0.28758887460831584   0.7933224189248625   0.8057192358344601   0.7296390740069862   0.016323775392647667   0.31182798955781615
0.07019072014605804   0.532827557517447   0.15179453717284652   0.028340211270525852   0.9036231039662386   0.9774802350592554   0.8068699122065681   0.4468777079216908   0.8087240948005411   0.9932349908929372   0.8072575185129988   0.37347203823500086   0.3066851719724417   0.4375123959860399   0.9627420225537898   0.04751378433632293   0.4676632477737703   0.6746157739860748   0.675153147945474   0.2541913654114604   0.6619440119393102   0.9449766999790885   0.6588293725528264   0.9423633758536443   0.5917532917932521   0.41214914246164147   0.5070348353799798   0.9140231645831184   0.6881301878270135   0.434668907402386   0.7001649231734116   0.46714545666142765   0.8794060930264724   0.4414339165094488   0.8929074046604129   0.09367341842642679   0.5727209210540307   0.003921520523408853   0.930165382106623   0.04615963409010386   0.10505767328026042   0.32930574653733413   0.25501223416114904   0.7919682686786435   0.44311366134095026   0.3843290465582457   0.5961828616083228   0.8496048928249992   0.8513603695476982   0.9721799040966043   0.08914802622834295   0.9355817282418807   0.16323018172068465   0.5375109966942182   0.3889831030549313   0.46843627158045303   0.2838240886942122   0.0960770801847694   0.4960756983945184   0.37476285315402624   0.7111031676401816   0.09215555966136055   0.5659103162878953   0.32860321906392237
0.6060454943599212   0.7628498131240264   0.3108980821267463   0.536634950385279   0.16293183301897082   0.3785207665657807   0.7147152205184236   0.6870300575602798   0.3115714634712726   0.4063408624691765   0.6255671942900806   0.7514483293183991   0.148341281750588   0.8688298657749584   0.2365840912351493   0.2830120577379461   0.8645171930563758   0.7727527855901889   0.7405083928406309   0.9082492045839199   0.15341402541619423   0.6805972259288283   0.17459807655273554   0.5796459855199975   0.5473685310562731   0.917747412804802   0.8636999944259892   0.0430110351347185   0.3844366980373023   0.5392266462390213   0.14898477390756565   0.3559809775744387   0.07286523456602965   0.13288578376984472   0.523417579617485   0.6045326482560396   0.9245239528154416   0.2640559179948864   0.28683348838233574   0.32152059051809345   0.0600067597590659   0.49130313240469753   0.5463250955417048   0.41327138593417356   0.9065927343428717   0.8107059064758692   0.3717270189889693   0.8336254004141761   0.35922420328659854   0.8929584936710672   0.5080270245629801   0.7906143652794576   0.9747875052492962   0.3537318474320459   0.3590422506554144   0.43463338770501897   0.9019222706832666   0.2208460636622012   0.8356246710379294   0.8301007394489794   0.9773983178678249   0.9567901456673148   0.5487911826555937   0.508580148930886
0.917391558108759   0.46548701326261727   0.0024660871138888277   0.0953087629967124   0.010798823765887353   0.6547811067867482   0.6307390681249195   0.26168336258253627   0.6515746204792888   0.761822613115681   0.12271204356193947   0.47106899730307866   0.6767871152299926   0.40809076568363506   0.763669792906525   0.03643560959805968   0.774864844546726   0.18724470202143387   0.9280451218685957   0.20633487014908025   0.797466526678901   0.23045455635411913   0.37925393921300204   0.6977547212181943   0.880074968570142   0.7649675430915018   0.3767878520991132   0.6024459582214818   0.8692761448042547   0.11018643630475372   0.7460487839741937   0.3407625956389456   0.2177015243249659   0.3483638231890728   0.6233367404122542   0.869693598335867   0.5409144090949733   0.9402730575054377   0.8596669475057291   0.8332579887378073   0.7660495645482474   0.7530283554840038   0.9316218256371335   0.6269231185887271   0.9685830378693463   0.5225737991298847   0.5523678864241314   0.9291683973705328   0.08850806929920423   0.7576062560383828   0.1755800343250182   0.32672243914905086   0.21923192449494952   0.6474198197336292   0.4295312503508245   0.9859598435101052   0.0015304001699836356   0.2990559965445564   0.8061945099385703   0.11626624517423828   0.46061599107501033   0.3587829390391187   0.9465275624328412   0.28300825643643096
0.6945664265267629   0.6057545835551149   0.014905736795707721   0.656085137847704   0.7259833886574167   0.08318078442523016   0.4625378503715763   0.7269167404771711   0.6374753193582124   0.3255745283868473   0.2869578160465581   0.4001943013281203   0.41824339486326295   0.6781547086532181   0.8574265656957336   0.41423445781801504   0.4167129946932793   0.3790987121086618   0.05123205575716324   0.29796821264377676   0.956097003618269   0.02031577306954313   0.10470449332432206   0.014959956207345785   0.261530577091506   0.4145611895144283   0.08979875652861434   0.35887481835964186   0.5355471884340893   0.3313804050891981   0.627260906157038   0.6319580778824707   0.8980718690758769   0.005805876702350793   0.34030309011047993   0.23176377655435038   0.4798284742126139   0.3276511680491326   0.4828765244147464   0.8175293187363354   0.06311547951933455   0.9485524559404708   0.43164446865758316   0.5195611060925586   0.10701847590106554   0.9282366828709276   0.3269399753332611   0.5046011498852128   0.8454878988095595   0.5136754933564994   0.23714121880464675   0.14572633152557096   0.30994071037547016   0.1822950882673013   0.6098803126476087   0.5137682536431003   0.41186884129959334   0.17648921156495048   0.2695772225371288   0.28200447708874987   0.9320403670869795   0.8488380435158179   0.7867006981223824   0.46447515835241454
0.868924887567645   0.900285587575347   0.35505622946479926   0.9449140522598559   0.7619064116665794   0.9720489047044194   0.028116254131538166   0.44031290237464316   0.9164185128570199   0.45837341134792003   0.7909750353268914   0.2945865708490722   0.6064778024815497   0.27607832308061875   0.18109472267928273   0.780818317205972   0.19460896118195634   0.09958911151566827   0.9115175001421539   0.498813840117222   0.2625685940949769   0.25075106799985036   0.12481680201977156   0.03433868176480746   0.39364370652733194   0.35046548042450326   0.7697605725549723   0.08942462950495152   0.6317372948607526   0.37841657572008386   0.7416443184234341   0.6491117271303084   0.7153187820037327   0.9200431643721638   0.9506692830965427   0.3545251562812362   0.10884097952218304   0.6439648412915451   0.76957456041726   0.5737068390752643   0.9142320183402267   0.5443757297758768   0.8580570602751061   0.07489299895804233   0.6516634242452498   0.29362466177602636   0.7332402582553345   0.04055431719323486   0.2580197177179179   0.9431591813515231   0.9634796857003621   0.9511296876882833   0.6262824228571653   0.5647426056314393   0.221835367276928   0.302017960557975   0.9109636408534325   0.6446994412592755   0.2711660841803853   0.9474928042767388   0.8021226613312495   0.0007345999677304108   0.5015915237631253   0.3737859652014744
0.8878906429910228   0.4563588701918536   0.6435344634880192   0.2988929662434321   0.23622721874577302   0.16273420841582725   0.9102942052326847   0.2583386490501972   0.9782075010278551   0.21957502706430415   0.9468145195323225   0.3072089613619139   0.3519250781706899   0.6548324214328649   0.7249791522553946   0.005191000803938933   0.44096143731725734   0.010132980173589433   0.4538130680750092   0.05769819652720021   0.6388387759860078   0.009398380205859022   0.952221544311884   0.6839122313257258   0.750948132994985   0.5530395100140054   0.30868708082386476   0.3850192650822937   0.5147209142492121   0.3903053015981781   0.39839287559118003   0.12668061603209652   0.5365134132213568   0.170730274533874   0.45157835605885743   0.8194716546701827   0.18458833505066696   0.5158978531010091   0.726599203803463   0.8142806538662437   0.7436268977334096   0.5057648729274197   0.2727861357284537   0.7565824573390435   0.10478812174740176   0.49636649272156064   0.32056459141656973   0.07267022601331768   0.35383998875241673   0.9433269827075552   0.011877510592705023   0.687650960931024   0.8391190745032047   0.5530216811093771   0.6134846350015251   0.5609703448989275   0.30260566128184785   0.38229140657550315   0.16190627894266757   0.7414986902287448   0.1180173262311809   0.866393553474494   0.43530707513920464   0.9272180363625011
0.37439042849777127   0.36062868054707437   0.1625209394107509   0.17063557902345763   0.2696023067503695   0.8642621878255137   0.8419563479941812   0.09796535301013994   0.9157623179979528   0.9209352051179585   0.8300788374014761   0.41031439207911596   0.07664324349474808   0.3679135240085813   0.2165942023999511   0.8493440471801885   0.7740375822129002   0.9856221174330781   0.054687923457283565   0.1078453569514437   0.6560202559817193   0.11922856395858414   0.6193808483180789   0.1806273205889426   0.28162982748394805   0.7585998834115097   0.456859908907328   0.009991741565484972   0.012027520733578507   0.8943376955859961   0.6149035609131469   0.912026388555345   0.09626520273562571   0.9734024904680376   0.7848247235116708   0.5017119964762291   0.01962195924087763   0.6054889664594564   0.5682305211117196   0.6523679492960406   0.24558437702797742   0.6198668490263782   0.513542597654436   0.5445225923445968   0.5895641210462581   0.5006382850677941   0.8941617493363571   0.3638952717556542   0.30793429356231006   0.7420384016562843   0.4373018404290291   0.35390353019016924   0.29590677282873157   0.8477007060702882   0.8223982795158822   0.4418771416348242   0.19964157009310582   0.8742982156022505   0.03757355600421148   0.9401651451585952   0.1800196108522282   0.2688092491427942   0.4693430348924919   0.28779719586255464
0.9344352338242508   0.648942400116416   0.9558004372380559   0.7432746035179578   0.3448711127779927   0.14830411504862195   0.061638687901698755   0.3793793317623036   0.03693681921568266   0.4062657133923377   0.6243368474726697   0.025475801572134325   0.7410300463869511   0.5585650073220495   0.8019385679567875   0.5835986599373101   0.5413884762938452   0.684266791719799   0.764365011952576   0.6434335147787149   0.3613688654416171   0.41545754257700473   0.29502197706008415   0.3556363189161603   0.4269336316173663   0.7665151424605887   0.3392215398220283   0.6123617153982025   0.0820625188393736   0.6182110274119668   0.27758285192032955   0.23298238363589893   0.04512569962369094   0.21194531401962907   0.6532460044476598   0.2075065820637646   0.3040956532367398   0.6533803066975796   0.8513074364908724   0.6239079221264545   0.7627071769428946   0.9691135149777806   0.08694242453829636   0.9804744073477395   0.40133831150127747   0.5536559724007759   0.7919204474782122   0.6248380884315793   0.9744046798839111   0.7871408299401871   0.4526989076561839   0.012476373033376719   0.8923421610445376   0.16892980252822035   0.17511605573585443   0.7794939893974778   0.8472164614208466   0.9569844885085913   0.5218700512881945   0.5719874073337132   0.5431208081841068   0.3036041818110117   0.6705626147973223   0.9480794852072587
0.7804136312412122   0.33449066683323103   0.5836201902590259   0.9676050778595191   0.3790753197399348   0.7808346944324552   0.7916997427808137   0.3427669894279399   0.4046706398560237   0.993693864492268   0.3390008351246297   0.3302906163945632   0.5123284788114861   0.8247640619640477   0.16388477938877527   0.5507966269970854   0.6651120173906395   0.8677795734554564   0.6420147281005807   0.9788092196633722   0.12199120920653274   0.5641753916444447   0.9714521133032584   0.03072973445611353   0.34157757796532046   0.2296847248112137   0.3878319230442326   0.0631246565965944   0.9625022582253857   0.44885003037875854   0.596132180263419   0.7203576671686545   0.557831618369362   0.45515616588649044   0.25713134513878927   0.3900670507740913   0.045503139557875855   0.6303921039224427   0.09324656575001401   0.8392704237770059   0.3803911221672363   0.7626125304669863   0.4512318376494333   0.8604612041136337   0.2583999129607036   0.19843713882254158   0.47977972434617483   0.8297314696575202   0.9168223349953831   0.9687524140113278   0.09194780130194223   0.7666068130609258   0.9543200767699974   0.5199023836325694   0.4958156210385233   0.046249145892271276   0.39648845840063546   0.0647462177460789   0.23868427589973398   0.6561820951181799   0.35098531884275963   0.43435411382363615   0.14543771014971996   0.816911671341174
0.9705941966755233   0.6717415833566498   0.6942058725002866   0.9564504672275403   0.7121942837148197   0.4733044445341083   0.21442614815411182   0.12671899757002014   0.7953719487194366   0.5045520305227804   0.12247834685216959   0.3601121845090944   0.8410518719494391   0.9846496468902111   0.6266627258136463   0.3138630386168231   0.44456341354880363   0.9199034291441321   0.38797844991391234   0.6576809434986431   0.09357809470604404   0.485549315320496   0.24254073976419238   0.8407692721574691   0.12298389803052075   0.8138077319638461   0.5483348672639057   0.8843188049299288   0.41078961431570105   0.3405032874297379   0.3339087191097939   0.7575998073599086   0.6154176655962644   0.8359512569069575   0.21143037225762434   0.39748762285081424   0.7743657936468253   0.8513016100167464   0.584767646443978   0.08362458423399116   0.3298023800980217   0.9313981808726143   0.19678919653006566   0.425943640735348   0.23622428539197765   0.4458488655521183   0.9542484567658732   0.585174368577879   0.11324038736145689   0.6320411335882721   0.40591358950196754   0.7008555636479502   0.7024507730457559   0.29153784615853423   0.07200487039217363   0.9432557562880415   0.08703310744949137   0.45558658925157675   0.8605744981345493   0.5457681334372273   0.31266731380266605   0.6042849792348304   0.2758068516905713   0.46214354920323614
0.9828649337046443   0.6728867983622161   0.07901765516050564   0.036199908467888106   0.7466406483126667   0.22703793281009782   0.12476919839463237   0.4510255398900092   0.6334002609512098   0.5949967992218257   0.7188556088926649   0.7501699762420591   0.930949487905454   0.30345895306329146   0.6468507385004912   0.8069142199540175   0.8439163804559626   0.8478723638117147   0.7862762403659419   0.2611460865167902   0.5312490666532965   0.24358738457688436   0.5104693886753706   0.7990025373135541   0.5483841329486522   0.5707005862146682   0.431451733514865   0.762802628845666   0.8017434846359855   0.3436626534045705   0.3066825351202326   0.3117770889556568   0.1683432236847757   0.7486658541827448   0.5878269262275678   0.5616071127135978   0.23739373577932174   0.44520690111945327   0.9409761877270766   0.7546928927595803   0.39347735532335915   0.5973345373077386   0.15469994736113465   0.49354680624279007   0.8622282886700626   0.3537471527308542   0.6442305586857641   0.6945442689292359   0.3138441557214104   0.7830465665161859   0.21277882517089908   0.93174164008357   0.5121006710854249   0.43938391311161545   0.9060962900506665   0.6199645511279132   0.3437574474006492   0.6907180589288707   0.31826936382309867   0.05835743841431545   0.10636371162132743   0.2455111578094174   0.37729317609602214   0.30366454565473516
0.7128863562979683   0.6481766205016789   0.22259322873488746   0.8101177394119451   0.8506580676279057   0.2944294677708246   0.5783626700491235   0.11557347048270916   0.5368139119064954   0.5113829012546387   0.3655838448782243   0.18383183039913917   0.024713240821070504   0.07199898814302327   0.4594875548275579   0.5638672792712259   0.6809557934204213   0.3812809292141526   0.14121819100445915   0.5055098408569105   0.5745920817990939   0.13576977140473517   0.763925014908437   0.20184529520217534   0.8617057255011256   0.4875931509030563   0.5413317861735496   0.3917275557902302   0.011047657873219888   0.19316368313223167   0.9629691161244261   0.27615408530752106   0.4742337459667245   0.681780781877593   0.5973852712462019   0.09232225490838186   0.449520505145654   0.6097817937345696   0.137897716418644   0.5284549756371559   0.7685647117252327   0.2285008645204171   0.9966795254141848   0.022945134780245388   0.19397262992613876   0.09273109311568192   0.2327545105057478   0.8210998395780701   0.33226690442501317   0.6051379422126256   0.6914227243321982   0.42937228378783987   0.3212192465517933   0.4119742590803939   0.728453608207772   0.1532181984803188   0.8469855005850687   0.730193477202801   0.13106833696157016   0.06089594357193696   0.3974649954394147   0.12041168346823132   0.9931706205429262   0.532440967934781
0.628900283714182   0.8919108189478142   0.9964910951287413   0.5094958331545356   0.43492765378804327   0.7991797258321324   0.7637365846229935   0.6883959935764656   0.10266074936303013   0.19404178361950672   0.07231386029079531   0.25902370978862577   0.7814415028112368   0.7820675245391128   0.3438602520830233   0.10580551130830693   0.9344560022261681   0.05187404733631179   0.21279191512145312   0.04490956773636997   0.5369910067867534   0.9314623638680805   0.21962129457852694   0.5124685998015889   0.9080907230725713   0.039551544920266225   0.2231301994497856   0.0029727666470532486   0.47316306928452806   0.2403718190881339   0.4593936148267921   0.3145767730705876   0.37050231992149796   0.046330035468627184   0.38707975453599675   0.05555306328196189   0.589060817110261   0.2642625109295144   0.043219502452973464   0.949747551973655   0.654604814884093   0.2123884635932026   0.8304275873315203   0.904837984237285   0.11761380809733955   0.2809260997251221   0.6108062927529934   0.3923693844356961   0.20952308502476819   0.24137455480485592   0.3876760933032078   0.3893966177886428   0.7363600157402401   0.0010027357167220103   0.9282824784764158   0.0748198447180552   0.36585769581874217   0.9546727002480948   0.541202723940419   0.019266781436093304   0.7767968787084811   0.6904101893185804   0.4979832214874455   0.06951922946243834
0.12219206382438814   0.4780217257253778   0.6675556341559251   0.16468124522515334   0.004578255727048598   0.19709562600025568   0.056749341402931745   0.7723118607894572   0.7950551707022804   0.9557210711953997   0.6690732480997239   0.3829152430008144   0.05869515496204027   0.9547183354786778   0.7407907696233081   0.3080953982827592   0.6928374591432981   0.00004563523058292627   0.1995880456828892   0.2888286168466659   0.916040580434817   0.3096354459120025   0.7016048241954437   0.21930938738422756   0.7938485166104289   0.8316137201866247   0.034049190039518513   0.05462814215907423   0.7892702608833803   0.6345180941863691   0.9772998486365868   0.282316281369617   0.9942150901810999   0.6787970229909692   0.30822660053686285   0.8994010383688026   0.9355199352190595   0.7240786875122915   0.5674358309135547   0.5913056400860434   0.24268247607576146   0.7240330522817086   0.3678477852306654   0.3024770232393775   0.3266418956409445   0.4143976063697061   0.6662429610352217   0.0831676358551499   0.5327933790305157   0.5827838861830814   0.6321937709957033   0.02853949369607567   0.7435231181471355   0.9482657919967123   0.6548939223591165   0.7462232123264587   0.7493080279660356   0.2694687690057431   0.3466673218222536   0.8468221739576561   0.813788092746976   0.5453900814934516   0.779231490908699   0.2555165338716127
0.5711056166712145   0.821357029211743   0.41138370567803356   0.9530395106322352   0.24446372103027006   0.406959422842037   0.7451407446428118   0.8698718747770854   0.7116703419997544   0.8241755366589556   0.11294697364710857   0.8413323810810097   0.968147223852619   0.8759097446622433   0.4580530512879921   0.09510916875455101   0.2188391958865834   0.6064409756565001   0.11138572946573846   0.24828699479689492   0.40505110313960735   0.06105089416304848   0.33215423855703946   0.9927704609252822   0.8339454864683928   0.23969386495130543   0.9207705328790059   0.03973095029304692   0.5894817654381227   0.8327344421092684   0.1756297882361941   0.16985907551596158   0.8778114234383684   0.008558905450312832   0.06268281458908553   0.32852669443495186   0.9096641995857494   0.1326491607880696   0.6046297633010934   0.23341752568040086   0.690825003699166   0.5262081851315695   0.493244033835355   0.985130530883506   0.2857739005595586   0.465157290968521   0.1610897952783155   0.9923600699582238   0.4518284140911658   0.22546342601721558   0.2403192623993096   0.9526291196651768   0.862346648653043   0.39272898390794714   0.06468947416311549   0.7827700441492152   0.9845352252146747   0.3841700784576343   0.002006659574029969   0.4542433497142634   0.07487102562892535   0.2515209176695647   0.39737689627293654   0.22082582403386253
0.3840460219297594   0.7253127325379952   0.9041328624375816   0.2356952931503566   0.09827212137020078   0.26015544156947423   0.743043067159266   0.2433352231921328   0.646443707279035   0.03469201555225862   0.5027238047599565   0.2907061035269559   0.784097058625992   0.6419630316443115   0.438034330596841   0.5079360593777407   0.7995618334113173   0.25779295318667717   0.43602767102281104   0.053692709663477244   0.7246908077823919   0.006272035517112438   0.038650774749874474   0.8328668856296148   0.3406447858526325   0.2809593029791172   0.1345179123122929   0.5971715924792581   0.24237266448243172   0.020803861409643007   0.39147484515302683   0.3538363692871253   0.5959289572033968   0.9861118458573844   0.8887510403930703   0.06313026576016939   0.8118318985774048   0.3441488142130729   0.45071670979622935   0.5551942063824288   0.012270065166087543   0.08635586102639577   0.014689038773418334   0.5015014967189515   0.28757925738369566   0.08008382550928332   0.9760382640235439   0.6686346110893368   0.9469344715310631   0.7991245225301661   0.841520351711251   0.07146301861007867   0.7045618070486314   0.7783206611205231   0.4500455065582241   0.7176266493229533   0.10863284984523466   0.7922088152631387   0.5612944661651538   0.654496383562784   0.2968009512678299   0.4480600010500658   0.11057775636892445   0.0993021771803552
0.2845308861017423   0.36170414002367   0.09588871759550611   0.5978006804614037   0.9969516287180467   0.28162031451438674   0.11985045357196225   0.9291660693720669   0.05001715718698355   0.4824957919842206   0.2783301018607113   0.8577030507619883   0.34545535013835216   0.7041751308636975   0.8282845953024871   0.1400764014390349   0.2368225002931175   0.9119663156005587   0.26699012913733333   0.485580017876251   0.9400215490252876   0.46390631455049297   0.1564123727684089   0.38627784069589577   0.6554906629235453   0.10220217452682295   0.0605236551729028   0.7884771602344921   0.6585390342054985   0.8205818600124363   0.9406732016009406   0.8593110908624252   0.608521877018515   0.3380860680282156   0.6623430997402292   0.0016080401004369392   0.26306652688016285   0.6339109371645181   0.8340585044377421   0.861531638661402   0.02624402658704539   0.7219446215639593   0.5670683753004088   0.37595162078515104   0.08622247756175778   0.2580383070134663   0.41065600253199985   0.9896737800892553   0.43073181463821253   0.15583613248664338   0.35013234735909704   0.20119661985476323   0.7721927804327139   0.33525427247420714   0.4094591457581565   0.34188552899233804   0.1636709034141989   0.9971682044459915   0.7471160460179272   0.3402774888919011   0.900604376534036   0.3632572672814734   0.9130575415801852   0.4787458502304991
0.8743603499469906   0.641312645717514   0.3459891662797764   0.10279422944534801   0.7881378723852328   0.3832743387040477   0.9353331637477765   0.11312044935609271   0.35740605774702033   0.22743820621740435   0.5852008163886795   0.9119238295013294   0.5852132773143064   0.8921839337431973   0.175741670630523   0.5700383005089914   0.42154237390010746   0.8950157292972057   0.4286256246125958   0.22976081161709033   0.5209379973660715   0.5317584620157324   0.5155680830324106   0.7510149613865913   0.6465776474190807   0.8904458162982183   0.16957891675263428   0.6482207319412433   0.8584397750338479   0.5071714775941706   0.23424575300485773   0.5351002825851505   0.5010337172868276   0.27973327137676623   0.6490449366161782   0.6231764530838211   0.9158204399725212   0.38754933763356897   0.4733032659856552   0.05313815257482963   0.4942780660724137   0.4925336083363632   0.044677641373059414   0.8233773409577393   0.9733400687063423   0.9607751463206309   0.5291095583406488   0.07236237957114805   0.32676242128726146   0.07032933002241258   0.35953064158801445   0.4241416476299048   0.4683226462534136   0.563157852428242   0.12528488858315673   0.8890413650447543   0.9672889289665859   0.2834245810514758   0.4762399519669785   0.2658649119609332   0.051468488994064775   0.8958752434179068   0.0029366859813232983   0.21272675938610355
0.5571904229216511   0.4033416350815436   0.9582590446082638   0.3893494184283643   0.5838503542153087   0.4425664887609127   0.4291494862676151   0.31698703885721624   0.25708793292804727   0.3722371587385001   0.06961884467960067   0.8928453912273114   0.7887652866746337   0.809079306310258   0.944333956096444   0.003804026182557169   0.8214763577080477   0.5256547252587823   0.46809400412946545   0.737939114221624   0.770007868713983   0.6297794818408755   0.46515731814814215   0.5252123548355204   0.21281744579233194   0.2264378467593319   0.5068982735398783   0.13586293640715613   0.6289670915770231   0.7838713579984192   0.07774878727226311   0.81887589754994   0.37187915864897586   0.4116341992599191   0.008129942592662446   0.9260305063226285   0.5831138719743422   0.602554892949661   0.06379598649621851   0.9222264801400714   0.7616375142662943   0.07690016769087873   0.5957019823667531   0.18428736591844735   0.9916296455523114   0.44712068585000325   0.13054466421861094   0.659075011082927   0.7788121997599794   0.22068283909067138   0.6236463906787327   0.5232120746757708   0.14984510818295627   0.43681148109225215   0.5458976034064695   0.7043361771258309   0.7779659495339803   0.025177281832333056   0.5377676608138071   0.7783056708032023   0.19485207755963826   0.42262238888267206   0.47397167431758863   0.856079190663131
0.4332145632933439   0.3457222211917933   0.8782696919508356   0.6717918247446837   0.44158491774103253   0.8986015353417901   0.7477250277322246   0.012716813661756733   0.6627727179810531   0.6779186962511187   0.12407863705349192   0.48950473898598595   0.5129276097980968   0.24110721515886652   0.5781810336470223   0.785168561860155   0.7349616602641165   0.21592993332653346   0.040413372833215236   0.006862891056952685   0.5401095827044782   0.7933075444438614   0.5664416985156266   0.15078370039382163   0.10689501941113429   0.4475853232520681   0.688172006564791   0.478991875649138   0.6653101016701017   0.548983787910278   0.9404469788325664   0.4662750619873812   0.0025373836890485914   0.8710650916591594   0.8163683417790746   0.9767703230013953   0.4896097738909517   0.6299578765002929   0.2381873081320522   0.19160176114124025   0.7546481136268353   0.4140279431737594   0.19777393529883694   0.18473887008428755   0.21453853092235706   0.6207203987298979   0.6313322367832104   0.033955169690465914   0.10764351151122277   0.17313507547782983   0.9431602302184192   0.5549632940413279   0.442333409841121   0.6241512875675518   0.0027132513858527784   0.08868823205394671   0.4397960261520725   0.7530861959083924   0.18634490960677824   0.1119179090525514   0.9501862522611207   0.12312831940809957   0.948157601474726   0.9203161479113111
0.19553813863428549   0.7091003762343402   0.7503836661758891   0.7355772778270236   0.9809996077119284   0.08837997750444224   0.11905142939267876   0.7016221081365577   0.8733560962007056   0.9152449020266124   0.17589119917425952   0.14665881409522974   0.43102268635958463   0.2910936144590606   0.17317794778840673   0.05797058204128304   0.9912266602075122   0.5380074185506682   0.9868330381816285   0.9460526729887316   0.04104040794639145   0.41487909914256865   0.038675436706902454   0.025736525077420472   0.8455022693121059   0.7057787229082284   0.28829177053101335   0.2901592472503969   0.8645026616001775   0.6173987454037863   0.1692403411383346   0.5885371391138392   0.9911465653994719   0.7021538433771738   0.9933491419640751   0.44187832501860946   0.5601238790398873   0.4110602289181132   0.8201711941756684   0.3839077429773264   0.5688972188323751   0.873052810367445   0.8333381559940398   0.43785506998859475   0.5278568108859836   0.4581737112248764   0.7946627192871374   0.4121185449111743   0.6823545415738776   0.752394988316648   0.5063709487561241   0.12195929766077743   0.8178518799737001   0.13499624291286175   0.33713060761778946   0.5334221585469382   0.8267053145742282   0.4328423995356879   0.34378146565371437   0.0915438335283288   0.266581435534341   0.021782170617574717   0.523610271478046   0.7076360905510024
0.6976842167019659   0.1487293602501297   0.6902721154840061   0.26978102056240766   0.1698274058159823   0.6905556490252533   0.8956093961968687   0.8576624756512333   0.4874728642421047   0.9381606607086054   0.38923844744074465   0.7357031779904559   0.6696209842684046   0.8031644177957437   0.05210783982295521   0.20228101944351767   0.8429156696941764   0.37032201826005573   0.7083263741692408   0.11073718591518888   0.5763342341598354   0.348539847642481   0.18471610269119487   0.4031010953641865   0.8786500174578695   0.1998104873923513   0.4944439872071888   0.13332007480177885   0.7088226116418872   0.509254838367098   0.5988345910103201   0.2756575991505455   0.2213497473997825   0.5710941776584926   0.20959614356957543   0.5399544211600895   0.5517287631313779   0.7679297598627489   0.1574883037466202   0.3376734017165719   0.7088130934372016   0.39760774160269324   0.4491619295773794   0.22693621580138298   0.13247885927736613   0.04906789396021222   0.26444582688618445   0.8238351204371965   0.25382884181949666   0.849257406567861   0.7700018396789957   0.6905150456354177   0.5450062301776095   0.34000256820076297   0.1711672486686756   0.4148574464848722   0.323656482777827   0.7689083905422703   0.9615711050991002   0.8749030253247826   0.7719277196464491   0.0009786306795214075   0.80408280135248   0.5372296236082108
0.06311462620924753   0.6033708890768282   0.3549208717751006   0.31029340780682774   0.9306357669318814   0.554302995116616   0.09047504488891615   0.48645828736963126   0.6768069251123847   0.705045588548755   0.32047320520992045   0.7959432417342136   0.13180069493477525   0.3650430203479921   0.14930595654124482   0.38108579524934133   0.8081442121569482   0.5961346298057217   0.18773485144214463   0.5061827699245587   0.03621649251049918   0.5951559991262003   0.38365205008966463   0.968953146316348   0.9731018663012516   0.9917851100493722   0.028731178314564034   0.6586597385095202   0.04246609936937026   0.4374821149327562   0.9382561334256478   0.17220145113988897   0.3656591742569855   0.7324365263840011   0.6177829282157274   0.3762582094056754   0.23385847932221027   0.36739350603600907   0.4684769716744826   0.9951724141563341   0.425714267165262   0.7712588762302873   0.28074212023233797   0.4889896442317753   0.3894977746547628   0.17610287710408698   0.8970900701426733   0.5200364979154274   0.4163959083535112   0.18431776705471484   0.8683588918281093   0.8613767594059072   0.37392980898414097   0.7468356521219587   0.9301027584024614   0.6891753082660181   0.008270634727155415   0.014399125737957503   0.312319830186734   0.3129170988603428   0.7744121554049451   0.6470056197019485   0.8438428585122514   0.31774468470400874
0.3486978882396831   0.8757467434716611   0.5631007382799134   0.8287550404722334   0.9592001135849203   0.6996438663675741   0.6660106681372401   0.30871854255680603   0.542804205231409   0.5153260993128593   0.7976517763091308   0.44734178315089884   0.16887439624726816   0.7684904471909006   0.8675490179066694   0.7581664748848806   0.16060376152011274   0.7540913214529432   0.5552291877199355   0.4452493760245379   0.3861916061151676   0.10708570175099473   0.7113863292076841   0.12750469132052916   0.03749371787548448   0.2313389582793336   0.1482855909277707   0.2987496508482958   0.0782936042905642   0.5316950919117595   0.48227492279053064   0.9900311082914898   0.5354893990591552   0.0163689925989001   0.6846231464813999   0.5426893251405909   0.36661500281188697   0.24787854540799942   0.8170741285747305   0.7845228502557102   0.20601124129177423   0.49378722395505625   0.2618449408547951   0.3392734742311723   0.8198196351766066   0.3867015222040615   0.550458611647111   0.21176878291064316   0.7823259173011221   0.15536256392472791   0.40217302071934036   0.9130191320623474   0.7040323130105579   0.6236674720129685   0.9198980979288097   0.9229880237708576   0.16854291395140283   0.6072984794140683   0.23527495144740984   0.3802986986302667   0.8019279111395159   0.359419934006069   0.41820082287267935   0.5957758483745565
0.5959166698477417   0.8656327100510127   0.15635588201788428   0.25650237414338417   0.776097034671135   0.4789311878469512   0.6058972703707732   0.04473359123274099   0.9937711173700129   0.3235686239222233   0.20372424965143293   0.1317144591703936   0.289738804359455   0.6999011519092548   0.2838261517226232   0.20872643539953598   0.12119589040805213   0.09260267249518643   0.04855120027521338   0.8284277367692693   0.31926797926853623   0.7331827384891174   0.630350377402534   0.23265188839471276   0.7233513094207946   0.8675500284381047   0.4739944953846497   0.9761495142513286   0.9472542747496595   0.3886188405911535   0.8680972250138764   0.9314159230185877   0.9534831573796466   0.06505021666893017   0.6643729753624436   0.799701463848194   0.6637443530201916   0.36514906475967535   0.3805468236398203   0.590975028448658   0.5425484626121395   0.2725463922644889   0.3319956233646069   0.7625472916793887   0.2232804833436033   0.5393636537753714   0.7016452459620729   0.529895403284676   0.49992917392280867   0.6718136253372667   0.22765075057742315   0.5537458890333474   0.5526748991731492   0.28319478474611326   0.3595535255635467   0.6223299660147598   0.5991917417935025   0.2181445680771831   0.6951805502011031   0.8226285021665658   0.9354473887733109   0.8529955033175077   0.31463372656128286   0.23165347371790773
0.39289892616117134   0.5804491110530188   0.982638103196676   0.46910618203851895   0.16961844281756808   0.04108545727764735   0.28099285723460304   0.939210778753843   0.6696892688947594   0.3692718319403806   0.05334210665717989   0.38546488972049553   0.11701436972161024   0.08607704719426731   0.6937885810936332   0.7631349237057358   0.5178226279281077   0.8679324791170842   0.99860803089253   0.94050642153917   0.5823752391547968   0.014936975799576445   0.6839743043312472   0.7088529478212623   0.18947631299362547   0.4344878647465576   0.7013362011345712   0.2397467657827433   0.019857870176057394   0.39340240746891025   0.4203433438999682   0.30053598702890033   0.350168601281298   0.02413057552852968   0.36700123724278827   0.9150710973084047   0.23315423155968776   0.9380535283342624   0.673212656149155   0.15193617360266903   0.7153316036315801   0.07012104921717817   0.674604625256625   0.21142975206349907   0.13295636447678325   0.05518407341760173   0.9906303209253778   0.5025768042422368   0.9434800514831577   0.6206962086710441   0.28929411979080666   0.26283003845949354   0.9236221813071004   0.22729380120213383   0.8689507758908385   0.9622940514305932   0.5734535800258024   0.20316322567360415   0.5019495386480501   0.04722295412218841   0.3402993484661146   0.2651096973393418   0.8287368824988951   0.8952867805195194
0.6249677448345345   0.1949886481221636   0.15413225724227003   0.6838570284560204   0.49201138035775127   0.1398045747045619   0.16350193631689214   0.1812802242137835   0.5485313288745935   0.5191083660335177   0.8742078165260855   0.9184501857542899   0.6249091475674932   0.29181456483138396   0.0052570406352470175   0.9561561343236967   0.05145556754169077   0.08865133915777977   0.5033075019871969   0.9089331802015084   0.7111562190755761   0.823541641818438   0.6745706194883018   0.013646399681988974   0.08618847424104163   0.6285529936962744   0.5204383622460318   0.3297893712259687   0.5941770938832903   0.4887484189917125   0.3569364259291396   0.14850914701218518   0.04564576500869682   0.9696400529581947   0.4827286094030541   0.2300589612578952   0.42073661744120366   0.6778254881268108   0.4774715687678071   0.27390282693419843   0.36928104989951294   0.589174148969031   0.9741640667806103   0.3649696467326901   0.6581248308239367   0.7656325071505931   0.29959344729230847   0.3513232470507011   0.5719363565828951   0.13707951345431865   0.7791550850462767   0.02153387582473247   0.9777592626996048   0.6483310944626062   0.42221865911713713   0.8730247288125473   0.9321134976909079   0.6786910415044114   0.939490049714083   0.6429657675546521   0.5113768802497043   0.0008655533776006526   0.46201848094627596   0.36906294062045364
0.14209583035019135   0.41169140440856966   0.48785441416566566   0.004093293887763541   0.4839709995262546   0.6460588972579766   0.1882609668733572   0.6527700468370624   0.9120346429433595   0.508979383803658   0.4091058818270804   0.63123617101233   0.9342753802437548   0.8606482893410519   0.9868872227099432   0.7582114421997826   0.0021618825528467943   0.1819572478366404   0.04739717299586024   0.11524567464513054   0.49078500230314254   0.18109169445903975   0.5853786920495843   0.7461827340246769   0.3486891719529512   0.7694002900504701   0.09752427788391861   0.7420894401369134   0.8647181724266966   0.12334139279249347   0.9092633110105615   0.08931939329985095   0.952683529483337   0.6143620089888355   0.5001574291834809   0.458083222287521   0.018408149239582304   0.7537137196477837   0.5132702064735377   0.6998717800877383   0.01624626668673551   0.5717564718111432   0.46587303347767745   0.5846261054426078   0.525461264383593   0.3906647773521035   0.8804943414280931   0.8384433714179309   0.17677209243064182   0.6212644873016334   0.7829700635441745   0.09635393128101759   0.3120539200039453   0.4979230945091399   0.8737067525336132   0.007034537981166645   0.3593703905206082   0.8835610855203044   0.37354932335013213   0.5489513156936456   0.3409622412810259   0.12984736587252077   0.8602791168765944   0.8490795356059073
0.3247159745942904   0.5580908940613776   0.394406083398917   0.2644534301632995   0.7992547102106974   0.16742611670927404   0.5139117419708238   0.4260100587453685   0.6224826177800556   0.5461616294076407   0.7309416784266493   0.3296561274643509   0.3104286977761103   0.04823853489850071   0.8572349258930361   0.3226215894831843   0.9510583072555021   0.16467744937819628   0.48368560254290394   0.7736702737895387   0.6100960659744762   0.03483008350567549   0.6234064856663095   0.9245907381836314   0.28538009138018583   0.47673918944429794   0.22900040226739254   0.6601373080203319   0.4861253811694884   0.30931307273502395   0.7150886602965688   0.2341272492749634   0.8636427633894328   0.7631514433273833   0.9841469818699196   0.9044711218106125   0.5532140656133224   0.7149129084288826   0.12691205597688343   0.5818495323274282   0.6021557583578203   0.5502354590506863   0.6432264534339794   0.8081792585378895   0.9920596923833441   0.5154053755450109   0.01981996776766996   0.8835885203542582   0.7066796010031583   0.03866618610071286   0.7908195655002774   0.22345121233392626   0.2205542198336699   0.729353113365689   0.07573090520370865   0.9893239630589629   0.3569114564442371   0.9662016700383056   0.09158392333378913   0.0848528412483504   0.8036973908309146   0.25128876160942304   0.9646718673569057   0.5030033089209223
0.20154163247309434   0.7010533025587368   0.32144541392292625   0.6948240503830326   0.20948194008975024   0.18564792701372593   0.30162544615525627   0.8112355300287745   0.502802339086592   0.14698174091301305   0.5108058806549789   0.5877843176948482   0.28224811925292204   0.4176286275473241   0.4350749754512702   0.5984603546358853   0.925336662808685   0.4514269575090185   0.3434910521174811   0.513607513387535   0.12163927197777027   0.20013819589959542   0.37881918476057536   0.01060420446661275   0.9200976395046759   0.4990848933408587   0.057373770837649156   0.31578015408358007   0.7106156994149256   0.31343696632713275   0.7557483246823928   0.5045446240548056   0.20781336032833375   0.1664552254141197   0.24494244402741402   0.9167603063599573   0.9255652410754117   0.7488265978667956   0.8098674685761438   0.318299951724072   0.00022857826672676362   0.2973996403577771   0.46637641645866273   0.804692438336537   0.8785893062889565   0.09726144445818166   0.08755723169808735   0.7940882338699242   0.9584916667842805   0.5981765511173229   0.030183460860438202   0.4783080797863442   0.24787596736935488   0.28473958479019024   0.2744351361780453   0.9737634557315387   0.04006260704102113   0.11828435937607053   0.029492692150631293   0.057003149371581276   0.11449736596560943   0.36945776150927495   0.21962522357448747   0.7387031976475092
0.11426878769888267   0.07205812115149787   0.7532488071158248   0.9340107593109723   0.23567948140992617   0.9747966766933163   0.6656915754177374   0.13992252544104802   0.2771878146256456   0.3766201255759932   0.6355081145572992   0.6616144456547038   0.029311847256290734   0.09188054078580303   0.3610729783792539   0.6878509899231653   0.9892492402152696   0.9735961814097325   0.33158028622862257   0.6308478405515839   0.8747518742496602   0.6041384199004576   0.1119550626541351   0.8921446429040747   0.7604830865507775   0.5320802987489597   0.35870625553831037   0.9581338835931024   0.5248036051408513   0.5572836220556434   0.693014680120573   0.8182113581520544   0.2476157905152057   0.1806634964796502   0.05750656556327378   0.1565969124973505   0.21830394325891497   0.08878295569384717   0.6964335871840199   0.46874592257418524   0.22905470304364536   0.11518677428411467   0.3648533009553973   0.8378980820226013   0.3543028287939852   0.5110483543836571   0.25289823830126223   0.9457534391185266   0.5938197422432077   0.9789680556346975   0.8941919827629519   0.9876195555254242   0.06901613710235639   0.42168443357905405   0.2011773026423789   0.1694081973733699   0.8214003465871507   0.24102093709940384   0.1436707370791051   0.012811284876019426   0.6030964033282358   0.15223798140555667   0.44723714989508523   0.5440653623018342
0.3740417002845904   0.037051207121442005   0.08238384893968788   0.7061672802792329   0.019738871490605162   0.5260028527377849   0.8294856106384256   0.7604138411607063   0.42591912924739744   0.5470347971030874   0.9352936278754738   0.772794285635282   0.35690299214504106   0.1253503635240334   0.7341163252330949   0.6033860882619121   0.5355026455578904   0.8843294264246295   0.5904455881539898   0.5905748033858926   0.9324062422296546   0.7320914450190729   0.14320843825890459   0.0465094410840585   0.5583645419450642   0.6950402378976309   0.06082458931921672   0.3403421608048256   0.5386256704544591   0.169037385159846   0.23133897868079106   0.5799283196441194   0.11270654120706165   0.6220025880567586   0.29604535080531724   0.8071340340088373   0.7558035490620206   0.49665222453272523   0.5619290255722224   0.20374794574692523   0.22030090350413023   0.6123227981080956   0.9714834374182325   0.6131731423610326   0.2878946612744756   0.8802313530890228   0.8282749991593279   0.5666637012769741   0.7295301193294114   0.1851911151913919   0.7674504098401113   0.22632154047214845   0.19090444887495223   0.016153730031545882   0.5361114311593201   0.6463932208280291   0.07819790766789056   0.3941511419747873   0.2400660803540029   0.8392591868191918   0.32239435860586996   0.8974989174420621   0.6781370547817805   0.6355112410722665
0.10209345510173971   0.2851761193339664   0.706653617363548   0.022338098711233993   0.8141987938272641   0.40494476624494363   0.87837861820422   0.45567439743425997   0.08466867449785279   0.21975365105355177   0.11092820836410885   0.22935285696211152   0.8937642256229006   0.2035999210220059   0.5748167772047887   0.5829596361340824   0.81556631795501   0.8094487790472186   0.3347506968507858   0.7437004493148907   0.49317195934914004   0.9119498616051566   0.6566136420690052   0.10818920824262412   0.3910785042474003   0.6267737422711901   0.9499600247054572   0.08585110953139014   0.5768797104201362   0.22182897602624643   0.07158140650123711   0.6301767120971302   0.49221103592228344   0.002075324972694661   0.9606531981371282   0.40082385513501867   0.5984468102993828   0.7984754039506887   0.38583642093233955   0.8178642190009362   0.7828804923443728   0.9890266249034702   0.051085724081553784   0.07416376968604559   0.2897085329952328   0.07707676329831367   0.3944720820125486   0.9659745614434214   0.8986300287478325   0.4503030210271236   0.44451205730709137   0.8801234519120313   0.32175031832769624   0.22847404500087715   0.37293065080585425   0.24994673981490115   0.8295392824054129   0.22639872002818248   0.412277452668726   0.8491228846798825   0.23109247210602996   0.42792331607749373   0.026441031736386452   0.03125866567894624
0.4482119797616571   0.4388966911740235   0.9753553076548327   0.9570948959929007   0.15850344676642428   0.3618199278757099   0.5808832256422841   0.9911203345494792   0.2598734180185918   0.9115169068485863   0.13637116833519272   0.11099688263744786   0.9381230996908956   0.6830428618477091   0.7634405175293384   0.8610501428225467   0.10858381728548273   0.4566441418195266   0.35116306486061244   0.011927258142664227   0.8774913451794528   0.028720825742032916   0.324722033124226   0.980668592463718   0.4292793654177957   0.5898241345680094   0.3493667254693933   0.02357369647081734   0.2707759186513714   0.2280042066922995   0.7684834998271092   0.03245336192133815   0.010902500632779599   0.3164872998437132   0.6321123314919165   0.9214564792838903   0.07277940094188405   0.6334444379960041   0.8686718139625781   0.06040633646134359   0.9641955836564013   0.17680029617647747   0.5175087491019656   0.04847907831867936   0.08670423847694853   0.14807947043444455   0.19278671597773966   0.06781048585496137   0.6574248730591529   0.5582553358664352   0.8434199905083464   0.04423678938414403   0.38664895440778146   0.3302511291741357   0.07493649068123714   0.01178342746280587   0.3757464537750018   0.013763829330422432   0.44282415918932067   0.09032694817891557   0.3029670528331178   0.38031939133441833   0.5741523452267426   0.02992061171757198
0.33877146917671647   0.20351909515794084   0.05664359612477694   0.9814415333988926   0.25206723069976794   0.05543962472349629   0.8638568801470373   0.9136310475439312   0.5946423576406151   0.4971842888570611   0.02043688963869092   0.8693942581597872   0.20799340323283366   0.16693315968292544   0.9455003989574537   0.8576108306969813   0.8322469494578318   0.15316933035250302   0.5026762397681331   0.7672838825180658   0.5292798966247141   0.7728499390180847   0.9285238945413905   0.7373632708004938   0.19050842744799756   0.5693308438601439   0.8718802984166136   0.7559217374016012   0.9384411967482296   0.5138912191366476   0.008023418269576338   0.84229068985767   0.3437988391076145   0.016706930279586436   0.9875865286308854   0.9728964316978828   0.13580543587478083   0.849773770596661   0.04208612967343164   0.11528560100090135   0.303558486416949   0.696604440244158   0.5394098899052985   0.34800171848283556   0.774278589792235   0.9237545012260733   0.610885995363908   0.6106384476823418   0.5837701623442374   0.35442365736592946   0.7390056969472943   0.8547167102807406   0.6453289655960078   0.8405324382292819   0.730982278677718   0.012426020423070673   0.3015301264883933   0.8238255079496954   0.7433957500468326   0.03952958872518797   0.16572469061361247   0.9740517373530345   0.7013096203734009   0.9242439877242866
0.8621662041966635   0.2774472971088765   0.16189973046810244   0.576242269241451   0.0878876144044285   0.3536927958828032   0.5510137351041945   0.9656038215591093   0.5041174520601911   0.9992691385168737   0.8120080381569001   0.11088711127836864   0.8587884864641833   0.15873670028759188   0.08102575947918217   0.09846109085529797   0.55725835997579   0.3349111923378964   0.3376300094323496   0.05893150213011001   0.3915336693621775   0.36085945498486194   0.6363203890589486   0.1346875144058234   0.529367465165514   0.08341215787598544   0.47442065859084626   0.5584452451643723   0.44147985076108553   0.7297193619931822   0.9234069234866518   0.5928414236052632   0.9373623987008944   0.7304502234763085   0.11139888532975158   0.48195431232689445   0.07857391223671117   0.5717135231887166   0.030373125850569414   0.3834932214715965   0.5213155522609212   0.2368023308508202   0.6927431164182198   0.3245617193414865   0.12978188289874368   0.8759428758659583   0.05642272735927116   0.1898742049356631   0.6004144177332297   0.7925307179899729   0.582002068768425   0.6314289597712908   0.15893456697214411   0.06281135599679061   0.6585951452817732   0.0385875361660276   0.22157216827124965   0.33236113252048216   0.5471962599520216   0.5566332238391332   0.14299825603453847   0.7606476093317656   0.5168231341014522   0.17314000236753666
0.6216827037736172   0.5238452784809453   0.8240800176832324   0.8485782830260502   0.4919008208748736   0.6479024026149871   0.7676572903239612   0.6587040780903871   0.891486403141644   0.8553716846250142   0.1856552215555363   0.02727511831909637   0.7325518361694998   0.7925603286282237   0.5270600762737631   0.9886875821530687   0.5109796678982502   0.4601991961077415   0.9798638163217415   0.4320543583139356   0.3679814118637117   0.699551586775976   0.4630406822202893   0.258914355946399   0.7462987080900945   0.17570630829503062   0.6389606645370569   0.4103360729203488   0.2543978872152209   0.5278039056800435   0.8713033742130957   0.7516319948299617   0.36291148407357693   0.6724322210550292   0.6856481526575594   0.7243568765108653   0.6303596479040772   0.8798718924268056   0.15858807638379632   0.7356692943577966   0.11937998000582693   0.41967269631906406   0.17872426006205483   0.303614936043861   0.7513985681421153   0.7201211095430881   0.7156835778417655   0.04470058009746198   0.0050998600520207596   0.5444148012480575   0.07672291330470861   0.6343645071771131   0.7507019728367998   0.016610895568013945   0.2054195390916129   0.8827325123471514   0.3877904887632229   0.3441786745129847   0.5197713864340535   0.1583756358362861   0.7574308408591458   0.4643067820861791   0.36118331005025717   0.4227063414784895
0.6380508608533189   0.04463408576711505   0.18245904998820234   0.11909140543462855   0.8866522927112036   0.32451297622402697   0.4667754721464368   0.07439082533716658   0.8815524326591829   0.7800981749759694   0.3900525588417282   0.4400263181600534   0.13085045982238303   0.7634872794079556   0.18463301975011528   0.557293805812902   0.7430599710591601   0.41930860489497085   0.6648616333160619   0.39891816997661583   0.9856291302000143   0.9550018228087918   0.30367832326580463   0.9762118284981264   0.3475782693466954   0.9103677370416767   0.12121927327760232   0.8571204230634978   0.46092597663549173   0.5858547608176498   0.6544438011311655   0.7827295977263312   0.5793735439763088   0.8057565858416802   0.26439124228943733   0.3427032795662778   0.44852308415392583   0.042269306433724695   0.07975822253932205   0.7854094737533759   0.7054631130947657   0.6229607015387538   0.4148965892232603   0.38649130377676   0.7198339828947514   0.6679588787299621   0.11121826595745561   0.4102794752786337   0.3722557135480561   0.7575911416882855   0.9899989926798533   0.5531590522151358   0.9113297369125644   0.17173638087063567   0.3355551915486878   0.7704294544888047   0.33195619293625545   0.36597979502895545   0.07116394925925044   0.4277261749225269   0.8834331087823296   0.32371048859523077   0.9914057267199284   0.6423167011691511
0.17796999568756386   0.700749787056477   0.5765091374966681   0.255825397392391   0.4581360127928124   0.032790908326514795   0.4652908715392125   0.8455459221137573   0.08588029924475632   0.27519976663822937   0.4752918788593592   0.2923868698986215   0.17455056233219202   0.1034633857675937   0.13973668731067146   0.5219574154098168   0.8425943693959366   0.7374835907386382   0.068572738051421   0.09423124048728991   0.959161260613607   0.4137731021434075   0.07716701133149262   0.45191453931813885   0.7811912649260431   0.7130233150869306   0.5006578738348245   0.19608914192574783   0.32305525213323066   0.6802324067604159   0.035367002295611974   0.35054321981199044   0.23717495288847434   0.4050326401221864   0.5600751234362528   0.05815634991336898   0.06262439055628234   0.30156925435459275   0.4203384361255813   0.5361989345035522   0.22003002116034578   0.5640856636159545   0.3517656980741603   0.4419676940162623   0.26086876054673885   0.15031256147254696   0.2745986867426677   0.9900531546981234   0.4796774956206958   0.43728924638561634   0.7739408129078432   0.7939640127723756   0.15662224348746515   0.7570568396252005   0.7385738106122313   0.4434207929603851   0.9194472905989908   0.3520241995030141   0.17849868717597844   0.3852644430470161   0.8568229000427084   0.05045494514842136   0.7581602510503972   0.849065508543464
0.6367928788823627   0.4863692815324669   0.40639455297623683   0.4070978145272017   0.3759241183356238   0.33605672005991993   0.13179586623356918   0.41704465982907823   0.8962466227149279   0.8987674736743035   0.357855053325726   0.6230806470567026   0.7396243792274628   0.14171063404910303   0.6192812427134947   0.17965985409631757   0.820177088628472   0.7896864345460889   0.44078255553751633   0.7943954110493014   0.9633541885857636   0.7392314893976676   0.6826223044871191   0.9453299025058375   0.32656130970340097   0.2528622078652007   0.2762277515108823   0.5382320879786358   0.9506371913677771   0.9168054878052808   0.14443188527731315   0.12118742814955755   0.054390568652849205   0.018038014130977224   0.7865768319515871   0.4981067810928549   0.31476618942538637   0.8763273800818742   0.1672955892380924   0.3184469269965373   0.4945891007969143   0.08664094553578527   0.7265130337005761   0.5240515159472359   0.5312349122111507   0.3474094561381177   0.04389072921345692   0.5787216134413984   0.2046736025077497   0.09454724827291702   0.7676629777025746   0.0404895254627626   0.25403641113997255   0.17774176046763623   0.6232310924252614   0.919302097313205   0.19964584248712333   0.159703746336659   0.8366542604736743   0.42119531622035017   0.884879653061737   0.2833763662547848   0.6693586712355819   0.10274838922381287
0.3902905522648227   0.19673542071899955   0.9428456375350058   0.578696873276577   0.859055640053672   0.8493259645808818   0.8989549083215489   0.9999752598351785   0.6543820375459223   0.7547787163079648   0.13129193061897426   0.959485734372416   0.40034562640594973   0.5770369558403285   0.5080608381937128   0.04018363705921093   0.2006997839188264   0.41733320950366953   0.6714065777200385   0.6189883208388608   0.31582013085708943   0.1339568432488847   0.0020479064844566683   0.5162399316150479   0.9255295785922668   0.9372214225298852   0.05920226894945088   0.9375430583384708   0.06647393853859478   0.08789545794900334   0.160247360627902   0.9375677985032923   0.4120919009926725   0.33311674164103855   0.028955430008927745   0.9780820641308763   0.011746274586722791   0.75607978580071   0.5208945918152149   0.9378984270716654   0.8110464906678964   0.33874657629704047   0.8494880140951764   0.31891010623280464   0.495226359810807   0.2047897330481558   0.8474401076107198   0.8026701746177568   0.5696967812185402   0.2675683105182706   0.7882378386612688   0.8651271162792858   0.5032228426799454   0.17967285256926727   0.6279904780333668   0.9275593177759935   0.09113094168727291   0.8465561109282287   0.5990350480244391   0.9494772536451173   0.07938466710055012   0.09047632512751871   0.07814045620922415   0.01157882657345186
0.26833817643265373   0.7517297488304783   0.22865244211404775   0.6926687203406472   0.7731118166218468   0.5469400157823224   0.38121233450332803   0.8899985457228904   0.20341503540330655   0.27937170526405186   0.5929744958420592   0.024871429443604553   0.7001921927233611   0.09969885269478458   0.9649840178086924   0.09731211166761097   0.6090612510360882   0.2531427417665559   0.36594896978425334   0.14783485802249371   0.5296765839355381   0.16266641663903716   0.2878085135750292   0.13625603144904186   0.26133840750288434   0.4109366678085589   0.0591560714609814   0.44358731110839467   0.4882265908810376   0.8639966520262364   0.6779437369576533   0.5535887653855042   0.28481155547773107   0.5846249467621846   0.08496924111559413   0.5287173359418996   0.58461936275437   0.48492609406740006   0.11998522330690174   0.4314052242742887   0.9755581117182818   0.23178335230084415   0.7540362535226485   0.283570366251795   0.44588152778274365   0.069116935661807   0.46622773994761924   0.1473143348027531   0.18454312027985928   0.6581802678532481   0.40707166848663784   0.7037270236943585   0.6963165293988217   0.7941836158270116   0.7291279315289845   0.15013825830885424   0.41150497392109064   0.20955866906482698   0.6441586904133904   0.6214209223669546   0.8268856111667207   0.724632574997427   0.5241734671064886   0.1900156980926659
0.8513274994484389   0.49284922269658277   0.7701372135838402   0.906445331840871   0.4054459716656953   0.4237322870347758   0.30390947363622095   0.7591309970381178   0.22090285138583599   0.7655520191815277   0.8968378051495831   0.055403973343759384   0.5245863219870143   0.9713684033545161   0.16770987362059858   0.9052657150349052   0.11308134806592368   0.7618097342896891   0.5235511832072082   0.28384479266795054   0.286195736899203   0.037177159292262195   0.9993777161007196   0.0938290945752846   0.4348682374507641   0.5443279365956795   0.22924050251687939   0.18738376273441365   0.029422265785068808   0.12059564956090364   0.9253310288806584   0.4282527656962958   0.8085194143992328   0.3550436303793759   0.02849322373107537   0.37284879235253643   0.28393309241221854   0.38367522702485984   0.8607833501104768   0.46758307731763127   0.17085174434629483   0.6218654927351707   0.33723216690326857   0.18373828464968076   0.8846560074470918   0.5846883334429085   0.337854450802549   0.08990919007439616   0.44978776999632775   0.04036039684722909   0.1086139482856696   0.9025254273399825   0.42036550421125896   0.9197647472863254   0.18328291940501115   0.4742726616436867   0.6118460898120262   0.5647211169069495   0.15478969567393577   0.1014238692911503   0.32791299739980756   0.18104588988208967   0.294006345563459   0.6338407919735191
0.15706125305351276   0.5591803971469189   0.9567741786601904   0.4501025073238383   0.27240524560642093   0.9744920637040104   0.6189197278576414   0.3601933172494421   0.8226174756100932   0.9341316668567814   0.5103057795719718   0.4576678899094596   0.4022519713988343   0.014366919570455917   0.32702286016696064   0.9833952282657729   0.7904058815868081   0.4496458026635064   0.17223316449302487   0.8819713589746225   0.4624928841870006   0.26859991278141676   0.8782268189295659   0.24813056700110356   0.3054316311334878   0.7094195156344978   0.9214526402693755   0.7980280596772653   0.03302638552706689   0.7349274519304874   0.3025329124117341   0.43783474242782316   0.2104089099169737   0.800795785073706   0.7922271328397622   0.9801668525183636   0.8081569385181394   0.7864288655032501   0.46520427267280157   0.9967716242525907   0.017751056931331253   0.33678306283974363   0.29297110817977673   0.11480026527796812   0.5552581727443306   0.06818315005832688   0.41474428925021084   0.8666696982768646   0.24982654161084286   0.3587636344238291   0.49329164898083533   0.06864163859959925   0.21680015608377595   0.6238361824933418   0.19075873656910128   0.6308068961717761   0.006391246166802273   0.8230403974196359   0.39853160372933905   0.6506400436534124   0.19823430764866284   0.03661153191638577   0.9333273310565374   0.6538684194008217
0.1804832507173316   0.6998284690766421   0.6403562228767608   0.5390681541228537   0.625225077973001   0.6316453190183152   0.2256119336265499   0.6723984558459891   0.3753985363621581   0.27288168459448614   0.7323202846457145   0.6037568172463899   0.1585983802783821   0.6490455021011444   0.5415615480766133   0.9729499210746138   0.15220713411157982   0.8260051046815086   0.14302994434727423   0.3223098774212013   0.953972826462917   0.7893935727651228   0.20970261329073678   0.6684414580203796   0.7734895757455854   0.08956510368848065   0.5693463904139761   0.12937330389752588   0.14826449777258446   0.4579197846701654   0.34373445678742615   0.45697484805153676   0.7728659614104264   0.18503810007567925   0.6114141721417116   0.8532180308051469   0.6142675811320443   0.5359925979745349   0.06985262406509833   0.8802681097305332   0.46206044702046445   0.7099874932930264   0.9268226797178241   0.5579582323093318   0.5080876205575474   0.9205939205279036   0.7171200664270874   0.8895167742889523   0.7345980448119621   0.8310288168394229   0.1477736760131113   0.7601434703914264   0.5863335470393777   0.37310903216925745   0.8040392192256851   0.3031686223398896   0.8134675856289513   0.18807093209357822   0.19262504708397357   0.44995059153474265   0.19920000449690695   0.6520783341190434   0.12277242301887523   0.5696824818042096
0.7371395574764426   0.942090840826017   0.1959497433010511   0.011724249494877704   0.22905193691889503   0.021496920298113488   0.47882967687396377   0.12220747520592544   0.49445389210693297   0.1904681034586906   0.33105600086085246   0.3620640048144991   0.9081203450675553   0.8173590712894332   0.5270167816351673   0.058895382474609466   0.09465275943860409   0.6292881391958549   0.33439173455119375   0.6089447909398669   0.8954527549416972   0.9772098050768115   0.21161931153231853   0.039262309135657286   0.15831319746525463   0.03511896425079457   0.015669568231267427   0.027538059640779586   0.9292612605463596   0.01362204395268108   0.5368398913573037   0.9053305844348541   0.43480736843942663   0.8231539404939905   0.20578389049645118   0.5432665796203551   0.5266870233718713   0.005794869204557319   0.6787671088612839   0.4843711971457456   0.4320342639332672   0.3765067300087024   0.34437537431009013   0.8754264062058789   0.5365815089915701   0.3992969249318908   0.13275606277777158   0.8361640970702215   0.37826831152631546   0.36417796068109626   0.11708649454650416   0.808626037429442   0.44900705097995586   0.35055591672841513   0.5802466031892005   0.9032954529945878   0.014199682540529229   0.5274019762344246   0.3744627126927493   0.36002887337423267   0.48751265916865794   0.5216071070298673   0.6956956038314654   0.8756576762284871
0.05547839523539071   0.145100377021165   0.3513202295213753   0.00023127002260825273   0.5188968862438206   0.7458034520892741   0.21856416674360374   0.16406717295238674   0.14062857471750517   0.3816254914081779   0.10147767219709958   0.35544113552294476   0.6916215237375493   0.031069574679762783   0.5212310690078991   0.452145682528357   0.6774218411970201   0.503667598445338   0.14676835631514978   0.0921168091541243   0.18990918202836216   0.9820604914154707   0.45107275248368434   0.21645913292563723   0.13443078679297146   0.8369601143943057   0.09975252296230903   0.21622786290302898   0.6155339005491508   0.09115666230503157   0.8811883562187053   0.05216068995064226   0.47490532583164563   0.7095311708968536   0.7797106840216057   0.6967195544276975   0.7832838020940963   0.6784615962170909   0.25847961501370664   0.24457387189934046   0.10586196089707627   0.17479399777175275   0.11171125869855686   0.15245706274521617   0.9159527788687141   0.19273350635628203   0.6606385062148725   0.935997929819579   0.7815219920757427   0.35577339196197627   0.5608859832525634   0.71977006691655   0.16598809152659183   0.2646167296569447   0.6796976270338582   0.6676093769659077   0.6910827656949462   0.5550855587600911   0.8999869430122525   0.9708898225382102   0.9077989636008499   0.8766239625430002   0.6415073279985458   0.7263159506388698
0.8019370027037735   0.7018299647712475   0.5297960692999889   0.5738588878936536   0.8859842238350595   0.5090964584149654   0.8691575630851164   0.6378609580740746   0.1044622317593168   0.15332306645298915   0.30827157983255293   0.9180908911575247   0.938474140232725   0.8887063367960445   0.6285739527986948   0.250481514191617   0.24739137453777882   0.33362077803595336   0.7285870097864423   0.27959169165340686   0.339592410936929   0.4569968154929531   0.0870796817878965   0.5532757410145371   0.5376554082331554   0.7551668507217056   0.5572836124879076   0.9794168531208836   0.6516711843980959   0.24607039230674016   0.6881260494027911   0.3415558950468089   0.5472089526387791   0.092747325853751   0.37985446957023816   0.42346500388928415   0.6087348124060541   0.20404098905770657   0.7512805167715434   0.17298348969766714   0.36134343786827533   0.8704202110217532   0.022693506985101076   0.8933917980442603   0.021751026931346357   0.4134233955288001   0.9356138251972046   0.3401160570297232   0.48409561869819095   0.6582565448070945   0.378330212709297   0.36069920390883964   0.832424434300095   0.4121861525003543   0.6902041633065059   0.019143308862030757   0.2852154816613159   0.3194388266466033   0.31034969373626775   0.5956783049727465   0.6764806692552617   0.11539783758889674   0.5590691769647244   0.42269481527507946
0.31513723138698646   0.24497762656714353   0.5363756699796233   0.5293030172308192   0.29338620445564007   0.8315542310383435   0.6007618447824187   0.18918696020109596   0.8092905857574492   0.17329768623124897   0.22243163207312167   0.8284877562922563   0.9768661514573541   0.7611115337308947   0.5322274687666158   0.8093444474302256   0.6916506697960382   0.44167270708429135   0.22187777503034803   0.21366614245747897   0.01517000054077643   0.3262748694953946   0.6628085980656238   0.7909713271823995   0.70003276915379   0.08129724292825105   0.12643292808600046   0.26166830995158036   0.4066465646981499   0.2497430118899076   0.5256710833035818   0.07248134975048441   0.5973559789407008   0.07644532565865866   0.3032394512304601   0.24399359345822808   0.6204898274833467   0.315333791927764   0.7710119824638443   0.43464914602800253   0.9288391576873085   0.8736610848434727   0.5491342074334963   0.22098300357052356   0.9136691571465321   0.5473862153480781   0.8863256093678726   0.43001167638812404   0.2136363879927421   0.466088972419827   0.7598926812818722   0.16834336643654366   0.8069898232945921   0.2163459605299194   0.23422159797829037   0.09586201668605925   0.20963384435389135   0.13990063487126073   0.9309821467478303   0.8518684232278312   0.5891440168705446   0.8245668429434967   0.15997016428398594   0.4172192771998286
0.6603048591832361   0.9509057581000241   0.6108359568504896   0.19623627362930507   0.746635702036704   0.40351954275194596   0.7245103474826171   0.7662245972411811   0.532999314043962   0.937430570332119   0.964617666200745   0.5978812308046374   0.7260094907493698   0.7210846098021996   0.7303960682224546   0.5020192141185782   0.5163756463954784   0.5811839749309388   0.7994139214746243   0.650150790890747   0.9272316295249338   0.7566171319874421   0.6394437571906383   0.23293151369091838   0.26692677034169765   0.805711373887418   0.028607800340148662   0.03669524006161331   0.5202910683049936   0.4021918311354721   0.3040974528575316   0.27047064282043226   0.9872917542610317   0.4647612608033531   0.33947978665678663   0.6725894120157948   0.26128226351166184   0.7436766510011535   0.6090837184343321   0.1705701978972167   0.7449066171161833   0.16249267607021475   0.8096697969597078   0.5204194070064697   0.8176749875912496   0.40587554408277265   0.17022603976906944   0.2874878933155513   0.5507482172495519   0.6001641701953546   0.14161823942892077   0.250792653253938   0.030457148944558317   0.19797233905988257   0.8375207865713892   0.9803220104335058   0.043165394683526676   0.7332110782565294   0.49804099991460254   0.3077325984177109   0.7818831311718648   0.9895344272553759   0.8889572814802705   0.1371624005204942
0.03697651405568146   0.8270417511851611   0.07928748452056275   0.6167429935140245   0.21930152646443188   0.4211662071023885   0.9090614447514933   0.32925510019847315   0.66855330921488   0.8210020369070339   0.7674432053225726   0.07846244694453515   0.6380961602703217   0.6230296978471512   0.9299224187511833   0.0981404365110294   0.5949307655867949   0.8898186195906218   0.43188141883658077   0.7904078380933185   0.8130476344149301   0.9002841923352459   0.5429241373563103   0.6532454375728243   0.7760711203592486   0.07324244115008478   0.4636366528357475   0.036502444058799835   0.5567695938948167   0.6520762340476963   0.5545752080842542   0.7072473438603266   0.8882162846799369   0.8310741971406624   0.7871320027616816   0.6287848969157915   0.2501201244096152   0.20804449929351115   0.8572095840104983   0.5306444604047621   0.6551893588228203   0.31822587970288935   0.4253281651739175   0.7402366223114436   0.8421417244078901   0.4179416873676434   0.8824040278176073   0.08699118473861928   0.0660706040486415   0.3446992462175586   0.4187673749818598   0.05048874067981944   0.5093010101538247   0.6926230121698623   0.8641921668976056   0.3432413968194928   0.6210847254738879   0.8615488150291999   0.07706016413592393   0.7144564999037013   0.3709646010642727   0.6535043157356887   0.21985058012542563   0.18381203949893918
0.7157752422414524   0.3352784360327994   0.7945224149515081   0.44357541718749555   0.8736335178335622   0.917336748665156   0.9121183871339008   0.3565842324488763   0.8075629137849208   0.5726375024475974   0.493351012152041   0.30609549176905687   0.29826190363109606   0.880014490277735   0.6291588452544354   0.9628540949495641   0.6771771781572082   0.018465675248535193   0.5520986811185116   0.2483975950458628   0.30621257709293553   0.3649613595128465   0.33224810099308594   0.06458555554692365   0.5904373348514831   0.029682923480047075   0.5377256860415778   0.6210101383594281   0.7168038170179207   0.11234617481489108   0.625607298907677   0.26442590591055176   0.909240903233   0.5397086723672937   0.13225628675563597   0.9583304141414949   0.6109789996019039   0.6596941820895587   0.5030974415012005   0.9954763191919308   0.9338018214446957   0.6412285068410234   0.9509987603826889   0.747078724146068   0.6275892443517602   0.2762671473281769   0.618750659389603   0.6824931685991443   0.03715190950027712   0.24658422384812986   0.08102497334802523   0.061483030239716276   0.32034809248235635   0.1342380490332388   0.4554176744403482   0.7970571243291645   0.41110718924935635   0.5945293766659451   0.32316138768471225   0.8387267101876695   0.8001281896474525   0.9348351945763865   0.8200639461835117   0.8432503909957387
0.8663263682027568   0.2936066877353631   0.8690651858008227   0.09617166684967073   0.23873712385099655   0.017339540407186133   0.2503145264112197   0.4136784982505264   0.2015852143507194   0.7707553165590563   0.16928955306319446   0.3521954680108101   0.8812371218683631   0.6365172675258175   0.7138718786228462   0.5551383436816456   0.4701299326190067   0.041987890859872354   0.390710490938134   0.7164116334939761   0.6700017429715542   0.10715269628348587   0.5706465447546223   0.8731612424982372   0.8036753747687976   0.8135460085481228   0.7015813589537995   0.7769895756485665   0.564938250917801   0.7962064681409367   0.4512668325425798   0.3633110773980402   0.3633530365670816   0.025451151581880382   0.28197727947938533   0.011115609387230082   0.4821159146987185   0.38893388405606294   0.5681054008565392   0.4559772657055845   0.011985982079711788   0.34694599319619057   0.17739490991840515   0.7395656322116084   0.3419842391081575   0.2397932969127047   0.6067483651637828   0.8664043897133712   0.53830886433936   0.4262472883645819   0.9051670062099834   0.08941481406480462   0.973370613421559   0.6300408202236453   0.4539001736674036   0.7261037366667644   0.6100175768544773   0.6045896686417649   0.1719228941880182   0.7149881272795343   0.1279016621557588   0.21565578458570198   0.603817493331479   0.25901086157394987
0.11591568007604701   0.8687097913895114   0.42642258341307393   0.5194452293623414   0.7739314409678895   0.6289164944768068   0.8196742182492911   0.6530408396489703   0.23562257662852956   0.2026692061122248   0.9145072120393076   0.5636260255841656   0.26225196320697064   0.5726283858885796   0.4606070383719041   0.8375222889174012   0.6522343863524933   0.9680387172468147   0.2886841441838859   0.12253416163786687   0.5243327241967345   0.7523829326611127   0.6848666508524068   0.863523300063917   0.4084170441206875   0.8836731412716012   0.25844406743933285   0.3440780707015756   0.634485603152798   0.25475664679479454   0.4387698491900418   0.6910372310526053   0.39886302652426847   0.052087440682569715   0.5242626371507341   0.12741120546843968   0.1366110633172978   0.4794590547939902   0.06365559877883001   0.2898889165510385   0.48437667696480446   0.5114203375471755   0.7749714545949441   0.1673547549131716   0.96004395276807   0.7590374048860629   0.09010480374253729   0.3038314548492546   0.5516269086473824   0.8753642636144616   0.8316607363032045   0.959753384147679   0.9171413054945844   0.6206076168196671   0.3928908871131626   0.2687161530950737   0.518278278970316   0.5685201761370975   0.8686282499624285   0.141304947626634   0.38166721565301814   0.08906112134310724   0.8049726511835985   0.8514160310755956
0.8972905386882137   0.5776407837959316   0.030001196588654386   0.684061276162424   0.9372465859201438   0.8186033789098688   0.939896392846117   0.38022982131316935   0.3856196772727613   0.9432391152954072   0.10823565654291266   0.4204764371654903   0.4684783717781769   0.32263149847573996   0.71534476942975   0.15176028407041667   0.950200092807861   0.7541113223386425   0.8467165194673215   0.010455336443782649   0.5685328771548428   0.6650502009955354   0.04174386828372303   0.1590393053681871   0.6712423384666292   0.0874094171996036   0.011742671695068645   0.47497802920576315   0.7339957525464854   0.2688060382897348   0.07184627884895156   0.09474820789259378   0.34837607527372405   0.32556692299432766   0.9636106223060389   0.6742717707271034   0.8798977034955472   0.0029354245185876857   0.24826585287628886   0.5225114866566868   0.9296976106876862   0.24882410217994513   0.4015493334089673   0.5120561502129041   0.36116473353284334   0.5837739011844099   0.3598054651252443   0.353016844844717   0.6899223950662142   0.4963644839848062   0.34806279343017565   0.8780388156389539   0.9559266425197288   0.22755844569507142   0.2762165145812241   0.7832906077463601   0.6075505672460046   0.9019915227007438   0.3126058922751852   0.10901883701925666   0.7276528637504576   0.899056098182156   0.06434003939889635   0.5865073503625698
0.7979552530627714   0.6502319960022109   0.662790705989929   0.07445120014966576   0.43679051952992803   0.06645809481780109   0.3029852408646847   0.7214343553049487   0.7468681244637139   0.5700936108329948   0.954922447434509   0.8433955396659949   0.7909414819439852   0.3425351651379234   0.678705932853285   0.06010493191963477   0.18339091469798044   0.4405436424371797   0.3661000405780997   0.9510860949003781   0.4557380509475229   0.5414875442550237   0.3017600011792034   0.3645787445378082   0.6577827978847515   0.8912555482528127   0.6389692951892744   0.2901275443881424   0.22099227835482346   0.8247974534350117   0.33598405432458966   0.5686931890831937   0.47412415389110957   0.2547038426020168   0.3810616068900806   0.7252976494171989   0.6831826719471245   0.9121686774640934   0.7023556740367957   0.665192717497564   0.49979175724914404   0.4716250350269136   0.33625563345869597   0.7141066225971859   0.04405370630162112   0.93013749077189   0.034495632279492615   0.34952787805937774   0.3862709084168696   0.038881942519077256   0.3955263370902182   0.059400333671235296   0.16527863006204616   0.21408448908406563   0.05954228276562857   0.4907071445880416   0.6911544761709366   0.9593806464820489   0.678480675875548   0.7654094951708428   0.00797180422381215   0.04721196901795556   0.9761250018387522   0.10021677767327869
0.5081800469746681   0.575586933991042   0.6398693683800563   0.38611015507609275   0.46412634067304703   0.645449443219152   0.6053737361005637   0.03658227701671499   0.0778554322561774   0.6065675007000747   0.20984739901034535   0.9771819433454797   0.9125768021941312   0.39248301161600907   0.1503051162447168   0.4864747987574381   0.22142232602319464   0.4331023651339602   0.4718244403691689   0.7210653035865954   0.21345052179938248   0.3858903961160047   0.49569943853041665   0.6208485259133166   0.7052704748247144   0.8103034621249627   0.8558300701503604   0.2347383708372239   0.24114413415166733   0.16485401890581072   0.25045633404979684   0.19815609382050892   0.16328870189548994   0.558286518205736   0.040608935039451455   0.22097415047502922   0.2507118997013587   0.16580350658972692   0.8903038187947346   0.7344993517175912   0.02928957367816408   0.7327011414557667   0.41847937842556576   0.013434048130995791   0.8158390518787816   0.346810745339762   0.9227799398951492   0.3925855222176792   0.11056857705406725   0.5365072832147993   0.06694986974478871   0.15784715138045524   0.8694244429024   0.3716532643089886   0.8164935356949918   0.9596910575599463   0.70613574100691   0.8133667461032525   0.7758846006555404   0.7387169070849171   0.4554238413055513   0.6475632395135257   0.8855807818608058   0.004217555367325956
0.4261342676273872   0.914862098057759   0.46710140343524   0.9907835072363301   0.6102952157486056   0.5680513527179969   0.5443214635400908   0.5981979850186511   0.4997266386945383   0.03154406950319758   0.47737159379530214   0.44035083363819577   0.6303021957921384   0.659890805194209   0.6608780581003103   0.48065977607824945   0.9241664547852284   0.8465240590909564   0.8849934574447699   0.7419428689933324   0.46874261347967716   0.1989608195774307   0.9994126755839641   0.7377253136260065   0.04260834585228996   0.28409872151967175   0.5323112721487241   0.7469418063896762   0.4323131301036844   0.7160473688016749   0.9879898086086332   0.14874382137102524   0.9325864914091461   0.6845032992984772   0.510618214813331   0.7083929877328294   0.3022842956170076   0.02461249410426827   0.8497401567130208   0.22773321165458   0.3781178408317792   0.1780884350133119   0.964746699268251   0.4857903426612476   0.909375227352102   0.9791276154358812   0.9653340236842869   0.7480650290352412   0.8667668814998121   0.6950288939162095   0.43302275153556286   0.0011232226455649109   0.4344537513961277   0.9789815251145346   0.44503294292692963   0.8523794012745397   0.5018672599869817   0.29447822581605737   0.9344147281135986   0.1439864135417102   0.19958296436997405   0.2698657317117891   0.08467457140057781   0.9162532018871302
0.8214651235381949   0.09177729669847721   0.11992787213232686   0.4304628592258826   0.9120898961860928   0.11264968126259603   0.15459384844803997   0.6823978301906415   0.04532301468628081   0.4176207873463866   0.7215710969124771   0.6812746075450765   0.6108692632901531   0.43863926223185196   0.2765381539855475   0.8288952062705368   0.10900200330317146   0.1441610364157946   0.34212342587194894   0.6849087927288267   0.9094190389331974   0.8742953047040055   0.2574488544713711   0.7686555908416964   0.08795391539500254   0.7825180080055283   0.13752098233904425   0.3381927316158138   0.17586401920890968   0.6698683267429323   0.9829271338910043   0.6557949014251724   0.13054100452262887   0.25224753939654565   0.2613560369785271   0.9745202938800959   0.5196717412324757   0.8136082771646936   0.9848178829929797   0.14562508760955903   0.4106697379293043   0.669447240748899   0.6426944571210307   0.46071629488073235   0.5012506989961069   0.7951519360448935   0.3852456026496596   0.692060704039036   0.41329678360110433   0.012633928039365298   0.24772462031061537   0.3538679724232221   0.23743276439219466   0.342765601296433   0.2647974864196111   0.6980730709980497   0.1068917598695658   0.09051806189988738   0.0034414494410839537   0.7235527771179538   0.5872200186370901   0.2769097847351937   0.018623566448104326   0.5779276895083948
0.17655028070778578   0.6074625439862946   0.37592910932707363   0.11721139462766242   0.6752995817116789   0.812310607941401   0.990683506677414   0.4251506905886265   0.2620027981105746   0.7996766799020357   0.7429588863667986   0.0712827181654044   0.024570033718379933   0.45691107860560265   0.47816139994718754   0.37320964716735466   0.9176782738488142   0.3663930167057153   0.4747199505061036   0.6496568700494009   0.33045825521172406   0.0894832319705216   0.4560963840579993   0.07172918054100606   0.15390797450393828   0.482020687984227   0.08016727473092566   0.9545177859133437   0.47860839279225936   0.669710080042826   0.08948376805351166   0.5293670953247172   0.21660559468168478   0.8700334001407902   0.346524881686713   0.45808437715931277   0.19203556096330485   0.4131223215351876   0.8683634817395255   0.08487472999195808   0.2743572871144907   0.046729304829472296   0.39364353123342183   0.4352178599425572   0.9438990319027666   0.9572460728589507   0.9375471471754225   0.36348867940155116   0.7899910573988284   0.4752253848747237   0.8573798724444969   0.4089708934882075   0.31138266460656894   0.8055153048318977   0.7678961043909852   0.8796037981634903   0.09477706992488417   0.9354819046911075   0.42137122270427224   0.42151942100417755   0.9027415089615793   0.5223595831559198   0.5530077409647468   0.3366446910122195
0.6283842218470886   0.47563027832644755   0.15936420973132492   0.9014268310696623   0.684485189944322   0.5183842054674969   0.22181706255590236   0.5379381516681112   0.8944941325454937   0.043158820592773164   0.36443719011140546   0.12896725817990365   0.5831114679389247   0.23764351576087547   0.5965410857204202   0.24936346001641332   0.48833439801404055   0.302161611069768   0.17516986301614804   0.8278440390122357   0.5855928890524612   0.7798020279138482   0.6221621220514012   0.49119934800001624   0.9572086672053726   0.3041717495874006   0.46279791232007633   0.5897725169303539   0.27272347726105056   0.7857875441199038   0.24098084976417397   0.05183436526224278   0.3782293447155569   0.7426287235271306   0.8765436596527685   0.9228671070823391   0.7951178767766323   0.5049852077662552   0.28000257393234823   0.6735036470659258   0.3067834787625917   0.20282359669648714   0.10483271091620022   0.8456596080536901   0.7211905897101305   0.42302156878263897   0.48267058886479897   0.35446026005367387   0.7639819225047579   0.11884981919523831   0.019872676544722634   0.7646877431233199   0.4912584452437073   0.33306227507533454   0.7788918267805487   0.7128533778610772   0.11302910052815042   0.5904335515482039   0.9023481671277802   0.789986270778738   0.3179112237515182   0.08544834378194871   0.6223455931954319   0.11648262371281218
0.011127744988926516   0.8826247470854616   0.5175128822792318   0.2708230156591221   0.28993715527879604   0.4596031783028226   0.03484229341443275   0.9163627556054482   0.5259552327740381   0.3407533591075843   0.014969616869710116   0.15167501248212836   0.034696787530330765   0.007691084032249815   0.23607779008916144   0.4388216346210512   0.9216676870021804   0.41725753248404596   0.33372962296138126   0.6488353638423132   0.6037564632506621   0.33180918870209725   0.7113840297659493   0.5323527401295011   0.5926287182617356   0.4491844416166356   0.1938711474867176   0.261529724470379   0.3026915629829396   0.989581263313813   0.15902885407228487   0.3451669688649307   0.7767363302089015   0.6488279042062287   0.14405923720257474   0.19349195638280234   0.7420395426785708   0.6411368201739789   0.9079814471134133   0.7546703217617511   0.8203718556763904   0.22387928768993295   0.574251824152032   0.10583495791943784   0.21661539242572825   0.8920700989878357   0.8628677943860827   0.5734822177899368   0.6239866741639927   0.44288565737120006   0.6689966468993651   0.3119524933195578   0.32129511118105303   0.45330439405738704   0.5099677928270803   0.9667855244546272   0.5445587809721515   0.8044764898511584   0.36590855562450547   0.7732935680718248   0.8025192382935807   0.1633396696771795   0.4579271085110922   0.018623246310073713
0.9821473826171904   0.9394603819872466   0.8836752843590602   0.9127882883906359   0.7655319901914621   0.04739028299941083   0.02080748997297743   0.3393060706006991   0.1415453160274695   0.6045046256282107   0.3518108430736123   0.027353577281141267   0.8202502048464164   0.15120023157082368   0.841843050246532   0.06056805282651413   0.27569142387426493   0.3467237417196653   0.47593449462202664   0.2872744847546893   0.47317218558068413   0.18338407204248583   0.018007386110934446   0.26865123844461564   0.49102480296349377   0.24392369005523928   0.1343321017518743   0.3558629500539797   0.7254928127720316   0.19653340705582845   0.11352461177889688   0.016556879453280656   0.5839474967445621   0.5920287814276177   0.7617137687052845   0.9892033021721394   0.7636972918981456   0.440828549856794   0.9198707184587525   0.9286352493456252   0.4880058680238807   0.09410480813712867   0.4439362238367258   0.6413607645909359   0.014833682443196545   0.9107207360946429   0.4259288377257914   0.3727095261463203   0.5238088794797028   0.6667970460394036   0.29159673597391705   0.016846576092340564   0.7983160667076712   0.4702636389835751   0.1780721241950202   0.0002896966390599099   0.21436856996310907   0.8782348575559574   0.41635835548973565   0.01108639446692052   0.45067127806496343   0.43740630769916344   0.4964876370309832   0.08245114512129527
0.9626654100410827   0.34330149956203476   0.0525514131942574   0.4410903805303593   0.9478317275978863   0.43258076346739194   0.626622575468466   0.06838085438403903   0.4240228481181834   0.7657837174279883   0.33502583949454895   0.05153427829169846   0.6257067814105123   0.29552007844441325   0.15695371529952878   0.05124458165263855   0.4113382114474031   0.4172852208884558   0.7405953598097932   0.04015818718571803   0.9606669333824397   0.9798789131892923   0.24410772277880993   0.9577070420644228   0.9980015233413569   0.6365774136272576   0.19155630958455255   0.5166166615340634   0.050169795743470705   0.20399665015986568   0.5649337341160865   0.4482358071500244   0.6261469476252873   0.43821293273187734   0.22990789462153755   0.39670152885832594   0.00044016621477504245   0.1426928542874641   0.07295417932200875   0.34545694720568737   0.5891019547673719   0.7254076333990083   0.3323588195122156   0.30529876001996936   0.6284350213849322   0.745528720209716   0.08825109673340566   0.3475917179555466   0.6304334980435753   0.10895130658245829   0.8966947871488531   0.8309750564214832   0.5802637023001046   0.9049546564225927   0.3317610530327666   0.38273924927145875   0.9541167546748173   0.46674172369071526   0.10185315841122905   0.9860377204131329   0.9536765884600422   0.32404886940325117   0.02889897908922031   0.6405807732074454
0.36457463369267035   0.5986412360042429   0.6965401595770047   0.3352820131874761   0.7361396123077382   0.8531125157945271   0.6082890628435991   0.9876902952319294   0.10570611426416288   0.7441612092120687   0.711594275694746   0.1567152388104463   0.5254424119640583   0.8392065527894762   0.37983322266197933   0.7739759895389875   0.571325657289241   0.3724648290987609   0.2779800642507503   0.7879382691258547   0.6176490688291988   0.04841595969550967   0.24908108516153   0.1473574959184093   0.2530744351365284   0.44977472369126675   0.5525409255845253   0.8120754827309332   0.5169348228287902   0.5966622078967397   0.9442518627409262   0.8243851874990038   0.41122870856462734   0.852500998684671   0.23265758704618025   0.6676699486885574   0.8857862966005691   0.013294445895194802   0.852824364384201   0.89369395914957   0.31446063931132806   0.6408296167964339   0.5748443001334506   0.10575569002371518   0.6968115704821293   0.5924136571009243   0.3257632149719206   0.9583981941053059   0.4437371353456009   0.14263893340965753   0.7732222893873953   0.1463227113743727   0.9268023125168107   0.5459767255129179   0.8289704266464691   0.32193752387536895   0.5155736039521833   0.6934757268282469   0.5963128396002889   0.6542675751868114   0.6297873073516143   0.6801812809330521   0.743488475216088   0.7605736160372416
0.31532666804028625   0.039351664136618135   0.16864417508263735   0.6548179260135264   0.6185150975581569   0.44693800703569386   0.8428809601107168   0.6964197319082205   0.17477796221255604   0.30429907362603636   0.0696586707233214   0.5500970205338478   0.24797564969574537   0.7583223481131185   0.24068824407685227   0.22815949665847887   0.732402045743562   0.06484662128487165   0.6443754044765634   0.5738919214716673   0.10261473839194775   0.3846653403518196   0.9008869292604754   0.8133183054344257   0.7872880703516615   0.3453136762152014   0.7322427541778381   0.1585003794208994   0.16877297279350456   0.8983756691795076   0.8893617940671213   0.4620806475126789   0.9939950105809485   0.5940765955534713   0.8197031233438   0.9119836269788311   0.7460193608852032   0.8357542474403526   0.5790148792669477   0.6838241303203522   0.013617315141641119   0.770907626155481   0.9346394747903843   0.10993220884868482   0.9110025767496934   0.3862422858036615   0.033752545529908855   0.29661390341425903   0.12371450639803187   0.04092860958846002   0.30150979135207073   0.13811352399335966   0.9549415336045274   0.14255294040895244   0.4121479972849494   0.6760328764806808   0.9609465230235789   0.5484763448554812   0.5924448739411494   0.7640492495018497   0.21492716213837568   0.7127220974151285   0.013429994674201676   0.08022511918149748
0.20130984699673454   0.9418144712596475   0.07879051988381737   0.9702929103328126   0.29030727024704117   0.555572185455986   0.04503797435390851   0.6736790069185536   0.1665927638490093   0.514643575867526   0.7435281830018378   0.535565482925194   0.21165123024448199   0.3720906354585735   0.3313801857168884   0.8595326064445132   0.25070470722090316   0.8236142906030923   0.738935311775739   0.09548335694266352   0.035777545082527486   0.1108921931879638   0.7255053171015373   0.015258237761166046   0.8344676980857929   0.16907772192831633   0.64671479721772   0.04496532742835339   0.5441604278387517   0.6135055364723303   0.6016768228638114   0.37128632050979976   0.37756766398974245   0.09886196060480433   0.8581486398619736   0.8357208375846058   0.16591643374526047   0.7267713251462308   0.5267684541450853   0.9761882311400926   0.9152117265243573   0.9031570345431384   0.7878331423693463   0.880704874197429   0.8794341814418298   0.7922648413551747   0.06232782526780898   0.865446636436263   0.04496648335603691   0.6231871194268583   0.41561302805008904   0.8204813090079096   0.5008060555172852   0.009681582954528038   0.8139362051862776   0.44919498849810985   0.1232383915275427   0.9108196223497237   0.9557875653243039   0.6134741509135041   0.9573219577822822   0.18404829720349292   0.4290191111792186   0.6372859197734114
0.042110231257924916   0.28089126266035447   0.6411859688098723   0.7565810455759824   0.16267604981609507   0.48862642130517975   0.5788581435420633   0.8911344091397194   0.11770956646005817   0.8654393018783214   0.16324511549197432   0.07065310013180977   0.616903510942773   0.8557577189237934   0.3493089103056967   0.6214581116336999   0.4936651194152303   0.9449380965740697   0.3935213449813928   0.007983960720195851   0.536343161632948   0.7608897993705768   0.9645022338021741   0.3706980409467844   0.49423293037502314   0.4799985367102223   0.32331626499230187   0.614116995370802   0.33155688055892807   0.9913721154050426   0.7444581214502385   0.7229825862310826   0.21384731409886992   0.12593281352672112   0.5812130059582642   0.6523294860992728   0.5969438031560969   0.27017509460292777   0.2319040956525675   0.030871374465572907   0.10327868374086659   0.3252369980288581   0.8383827506711747   0.022887413745377058   0.5669355221079185   0.5643471986582813   0.8738805168690005   0.6521893727985927   0.07270259173289535   0.08434866194805904   0.5505642518766987   0.0380723774277907   0.7411457111739673   0.0929765465430165   0.8061061304264601   0.3150897911967081   0.5272983970750974   0.9670437330162954   0.22489312446819584   0.6627603050974353   0.9303545939190004   0.6968686384133677   0.9929890288156283   0.6318889306318624
0.8270759101781339   0.3716316403845095   0.15460627814445366   0.6090015168864853   0.26014038807021533   0.8072844417262282   0.2807257612754532   0.9568121440878926   0.18743779633732   0.7229357797781691   0.7301615093987546   0.9187397666601019   0.4462920851633527   0.6299592332351527   0.9240553789722945   0.6036499754633938   0.9189936880882553   0.6629155002188573   0.6991622545040986   0.9408896703659585   0.9886390941692549   0.9660468618054896   0.7061732256884703   0.30900073973409614   0.16156318399112105   0.5944152214209801   0.5515669475440166   0.6999992228476108   0.9014227959209057   0.7871307796947519   0.27084118626856346   0.7431870787597181   0.7139849995835857   0.06419499991658276   0.5406796768698089   0.8244473120996162   0.267692914420233   0.4342357666814301   0.6166242978975144   0.22079733663622236   0.34869922633197764   0.7713202664625729   0.9174620433934157   0.2799076662702638   0.3600601321627227   0.8052734046570832   0.21128881770494554   0.9709069265361676   0.19849694817160168   0.2108581832361031   0.659721870160929   0.2709077036885568   0.297074152250696   0.4237274035413512   0.3888806838923655   0.5277206249288386   0.5830891526671103   0.35953240362476846   0.8482010070225566   0.7032733128292225   0.31539623824687724   0.9252966369433383   0.2315767091250422   0.48247597619300014
0.9666970119148997   0.15397637048076546   0.3141146657316264   0.20256830992273633   0.606636879752177   0.34870296582368226   0.10282584802668085   0.2316613833865687   0.4081399315805752   0.13784478258757912   0.4431039778657519   0.9607536796980118   0.11106577932987924   0.714117379046228   0.054223293973386426   0.43303305476917314   0.527976626662769   0.3545849754214595   0.20602228695082983   0.7297597419399506   0.21258038841589172   0.4292883384781212   0.9744455778257877   0.2472837657469505   0.2458833765009921   0.2753119679973557   0.6603309120941613   0.044715455824214136   0.6392464967488152   0.9266090021736735   0.5575050640674803   0.8130540724376455   0.23110656516824   0.7887642195860943   0.11440108620172847   0.8523003927396336   0.12004078583836075   0.07464684053986641   0.06017779222834205   0.4192673379704605   0.5920641591755917   0.7200618651184069   0.8541555052775123   0.6895075960305098   0.3794837707597   0.2907735266402857   0.8797099274517246   0.4422238302835594   0.13360039425870796   0.015461558642930015   0.21937901535756335   0.3975083744593452   0.4943538975098927   0.08885255646925655   0.661873951290083   0.5844543020216998   0.26324733234165276   0.3000883368831622   0.5474728650883545   0.7321539092820661   0.143206546503292   0.2254414963432958   0.48729507286001245   0.3128865713116057
0.5511423873277003   0.5053796312248889   0.6331395675825002   0.6233789752810959   0.1716586165680002   0.2146061045846032   0.7534296401307756   0.18115514499753646   0.038058222309292254   0.19914454594167316   0.5340506247732123   0.7836467705381912   0.5437043247993996   0.11029198947241661   0.8721766734831293   0.19919246851649144   0.28045699245774675   0.8102036525892544   0.3247038083947748   0.4670385592344253   0.13725044595445474   0.5847621562459586   0.8374087355347624   0.15415198792281962   0.5861080586267545   0.07938252502106968   0.2042691679522622   0.5307730126417238   0.4144494420587543   0.8647764204364665   0.45083952782148656   0.34961786764418734   0.37639121974946205   0.6656318744947933   0.9167889030482743   0.5659710971059961   0.8326868949500625   0.5553398850223767   0.04461222956514498   0.36677862858950466   0.5522299024923157   0.7451362324331223   0.7199084211703701   0.8997400693550793   0.41497945653786106   0.16037407618716373   0.8824996856356078   0.7455880814322597   0.8288713979111065   0.08099155116609405   0.6782305176833456   0.21481506879053597   0.41442195585235225   0.21621513072962756   0.22739098986185902   0.8651972011463487   0.03803073610289018   0.5505832562348342   0.3106020868135847   0.29922610404035255   0.20534384115282764   0.9952433712124574   0.2659898572484397   0.9324474754508478
0.6531139386605118   0.25010713877933516   0.5460814360780696   0.03270740609576848   0.23813448212265081   0.08973306259217143   0.6635817504424618   0.2871193246635087   0.4092630842115443   0.008741511426077367   0.9853512327591162   0.07230425587297273   0.994841128359192   0.7925263806964499   0.7579602428972572   0.20710705472662408   0.9568103922563018   0.24194312446161562   0.4473581560836725   0.9078809506862715   0.7514665511034743   0.24669975324915813   0.18136829883523276   0.9754334752354237   0.09835261244296238   0.996592614469823   0.6352868627571632   0.9427260691396552   0.8602181303203116   0.9068595518776515   0.9717051123147014   0.6556067444761465   0.4509550461087673   0.8981180404515742   0.9863538795555852   0.5833024886031738   0.4561139177495752   0.10559165975512438   0.22839363665832793   0.3761954338765497   0.49930352549327334   0.8636485352935087   0.7810354805746554   0.46831448319027813   0.7478369743897991   0.6169487820443507   0.5996671817394227   0.4928810079548544   0.6494843619468368   0.6203561675745276   0.9643803189822595   0.5501549388151992   0.7892662316265252   0.7134966156968761   0.9926752066675582   0.8945481943390527   0.3383111855177579   0.8153785752453019   0.006321327111972968   0.31124570573587895   0.8821972677681826   0.7097869154901775   0.7779276904536451   0.9350502718593292
0.3828937422749093   0.8461383801966688   0.9968922098789896   0.46673578866905113   0.6350567678851102   0.22918959815231812   0.39722502813956695   0.9738547807141967   0.9855724059382734   0.6088334305777905   0.43284470915730744   0.4236998418989975   0.19630617431174824   0.8953368148809144   0.44016950248974934   0.5291516475599448   0.8579949887939904   0.0799582396356125   0.43384817537777637   0.21790594182406586   0.9757977210258076   0.37017132414543497   0.6559204849241314   0.2828556699647366   0.5929039787508984   0.5240329439487662   0.6590282750451417   0.8161198812956855   0.9578472108657882   0.2948433457964481   0.26180324690557477   0.8422651005814887   0.9722748049275147   0.6860099152186576   0.8289585377482673   0.4185652586824912   0.7759686306157665   0.7906731003377433   0.388789035258518   0.8894136111225465   0.9179736418217762   0.7107148607021307   0.9549408598807416   0.6715076692984806   0.9421759207959685   0.3405435365566958   0.29902037495661027   0.38865199933374395   0.3492719420450701   0.8165105926079296   0.6399920999114685   0.5725321180380585   0.3914247311792819   0.5216672468114815   0.3781888530058937   0.7302670174565697   0.4191499262517671   0.8356573315928237   0.5492303152576264   0.3117017587740785   0.6431812956360006   0.04498423125508053   0.16044127999910843   0.4222881476515321
0.7252076538142245   0.33426937055294975   0.20550042011836683   0.7507804783530515   0.783031733018256   0.993725833996254   0.9064800451617566   0.3621284790193076   0.4337597909731859   0.17721524138832445   0.26648794525028807   0.7895963609812491   0.042335059793903985   0.655547994576843   0.8882990922443943   0.05932934352467933   0.6231851335421369   0.8198906629840192   0.3390687769867679   0.7476275847506008   0.9800038379061362   0.7749064317289387   0.17862749698765948   0.3253394370990687   0.25479618409191174   0.44063706117598894   0.9731270768692927   0.5745589587460171   0.4717644510736558   0.4469112271797349   0.06664703170753608   0.21243047972670953   0.03800466010046988   0.26969598579141046   0.800159086457248   0.42283411874546045   0.9956696003065659   0.6141479912145674   0.9118599942128537   0.3635047752207811   0.37248446676442903   0.7942573282305482   0.5727912172260857   0.6158771904701803   0.3924806288582928   0.019350896501609528   0.3941637202384263   0.29053775337111165   0.1376844447663811   0.5787138353256206   0.4210366433691336   0.7159787946250945   0.6659199936927254   0.13180260814588568   0.35438961166159755   0.503548314898385   0.6279153335922555   0.8621066223544752   0.5542305252043496   0.08071419615292454   0.6322457332856896   0.24795863113990774   0.6423705309914959   0.7172094209321435
0.2597612665212605   0.4537013029093595   0.06957931376541007   0.10133223046196309   0.8672806376629677   0.43435040640774997   0.6754155935269838   0.8107944770908514   0.7295961928965866   0.8556365710821294   0.25437895015785017   0.09481568246575693   0.06367619920386125   0.7238339629362437   0.8999893384962526   0.591267367567372   0.4357608656116058   0.8617273405817685   0.3457588132919031   0.5105531714144474   0.8035151323259162   0.6137687094418608   0.7033882823004073   0.793343750482304   0.5437538658046558   0.16006740653250123   0.6338089685349972   0.6920115200203409   0.6764732281416881   0.7257170001247513   0.9583933750080134   0.8812170429294894   0.9468770352451015   0.8700804290426218   0.7040144248501632   0.7864013604637325   0.8832008360412402   0.14624646610637818   0.8040250863539106   0.19513399289636058   0.4474399704296344   0.2845191255246097   0.4582662730620074   0.6845808214819131   0.6439248381037181   0.6707504160827489   0.7548779907616001   0.8912370709996091   0.10017097229906244   0.5106830095502477   0.12106902222660294   0.19922555097926822   0.4236977441573744   0.7849660094254964   0.16267564721858957   0.31800850804977876   0.47682070891227285   0.9148855803828745   0.4586612223684264   0.5316071475860462   0.5936198728710326   0.7686391142764963   0.6546361360145158   0.33647315468968564
0.1461799024413982   0.48411998875188667   0.19636986295250838   0.6518923332077725   0.50225506433768   0.8133695726691378   0.44149187219090824   0.7606552622081634   0.40208409203861756   0.30268656311889014   0.32042284996430526   0.5614297112288951   0.9783863478812432   0.5177205536933938   0.15774720274571571   0.24342120317911634   0.5015656389689703   0.6028349733105192   0.6990859803772894   0.7118140555930701   0.9079457660979378   0.8341958590340228   0.044449844362773556   0.37534090090338446   0.7617658636565395   0.35007587028213616   0.8480799814102652   0.7234485676956119   0.2595107993188595   0.5367062976129984   0.40658810921935695   0.9627933054874486   0.857426707280242   0.23401973449410826   0.08616525925505168   0.40136359425855345   0.8790403593989987   0.7162991808007145   0.928418056509336   0.1579423910794371   0.37747472043002833   0.11346420749019533   0.2293320761320466   0.446128335486367   0.46952895433209063   0.2792683484561725   0.18488223176927304   0.07078743458298256   0.7077630906755511   0.9291924781740363   0.33680225035900785   0.34733886688737065   0.4482522913566916   0.39248618056103796   0.9302141411396508   0.384545561399922   0.5908255840764497   0.1584664460669297   0.8440488818845993   0.9831819671413686   0.711785224677451   0.4421672652662152   0.9156308253752633   0.8252395760619314
0.3343105042474226   0.3287030577760198   0.6862987492432167   0.37911124057556445   0.864781549915332   0.049434709319847364   0.5014165174739437   0.30832380599258186   0.15701845923978083   0.12024223114581105   0.1646142671149358   0.9609849391052112   0.7087661678830892   0.7277560505847731   0.2344001259752849   0.5764393777052892   0.11794058380663963   0.5692896045178434   0.39035124409068567   0.5932574105639207   0.4061553591291887   0.12712233925162825   0.4747204187154224   0.7680178345019891   0.07184485488176613   0.7984192814756084   0.7884216694722057   0.38890659392642474   0.2070633049664342   0.7489845721557611   0.2870051519982621   0.08058278793384287   0.05004484572665335   0.62874234100995   0.12239088488332633   0.11959784882863161   0.3412786778435641   0.9009862904251769   0.8879907589080415   0.5431584711233424   0.22333809403692445   0.3316966859073335   0.4976395148173558   0.9499010605594218   0.8171827349077357   0.2045743466557052   0.022919096101933375   0.1818832260574326   0.7453378800259696   0.4061550651800968   0.23449742662972764   0.7929766321310079   0.5382745750595355   0.6571704930243357   0.9474922746314656   0.712393844197165   0.48822972933288206   0.02842815201438576   0.8251013897481392   0.5927959953685333   0.14695105148931797   0.12744186158920887   0.9371106308400977   0.04963752424519098
0.9236129574523936   0.7957451756818754   0.43947111602274197   0.0997364636857692   0.10643022254465777   0.5911708290261702   0.4165520199208086   0.9178532376283366   0.36109234251868816   0.1850157638460734   0.18205459329108095   0.12487660549732874   0.8228177674591527   0.5278452708217376   0.23456231865961544   0.41248276130016376   0.33458803812627064   0.4994171188073519   0.40946092891147623   0.8196867659316304   0.18763698663695266   0.371975257218143   0.4723502980713785   0.7700492416864394   0.26402402918455914   0.5762300815362676   0.03287918204863657   0.6703127780006701   0.15759380663990136   0.9850592525100974   0.616327162127828   0.7524595403723335   0.7965014641212133   0.800043488664024   0.43427256883674703   0.6275829348750048   0.9736836966620604   0.27219821784228637   0.19971025017713162   0.2151001735748411   0.6390956585357899   0.7727810990349345   0.7902493212656554   0.39541340764321076   0.45145867189883715   0.40080584181679146   0.3178990231942769   0.6253641659567714   0.18743464271427804   0.8245757602805239   0.28501984114564033   0.9550513879561012   0.02984083607437666   0.8395165077704265   0.6686926790178123   0.20259184758376764   0.23333937195316345   0.03947301910640249   0.23442011018106526   0.5750089127087628   0.25965567529110295   0.7672748012641162   0.03470986000393363   0.35990873913392174
0.6205600167553131   0.9944937022291817   0.24446053873827825   0.964495331490711   0.16910134485647596   0.5936878604123902   0.9265615155440013   0.3391311655339396   0.981666702142198   0.7691121001318663   0.6415416743983611   0.3840797775778384   0.9518258660678213   0.9295955923614398   0.9728489953805488   0.1814879299940708   0.7184864941146578   0.8901225732550373   0.7384288851994835   0.606479017285308   0.45883081882355486   0.12284777199092119   0.7037190251955499   0.24657027815138624   0.8382708020682418   0.12835406976173952   0.45925848645727163   0.2820749466606753   0.6691694572117658   0.5346662093493494   0.5326969709132703   0.9429437811267356   0.6875027550695678   0.765554109217483   0.8911552965149092   0.5588640035488972   0.7356768890017465   0.8359585168560433   0.9183063011343604   0.37737607355482644   0.017190394887088775   0.9458359436010059   0.1798774159348769   0.7708970562695184   0.5583595760635339   0.8229881716100848   0.47615839073932703   0.5243267781181322   0.7200887739952921   0.6946341018483452   0.01689990428205544   0.24225183145745696   0.05091931678352635   0.15996789249899585   0.48420293336878517   0.2993080503307213   0.3634165617139585   0.3944137832815128   0.5930476368538761   0.7404440467818241   0.6277396727122119   0.5584552664254696   0.6747413357195156   0.36306797322699763
0.6105492778251231   0.6126193228244636   0.4948639197846387   0.5921709169574791   0.05218970176158919   0.789631151214379   0.01870552904531162   0.0678441388393469   0.33210092776629707   0.09499704936603376   0.0018056247632561796   0.8255923073818899   0.28118161098277067   0.9350291568670379   0.517602691394471   0.5262842570511687   0.9177650492688122   0.5406153735855251   0.924555054540595   0.7858402102693446   0.2900253765566003   0.9821601071600555   0.24981371882107936   0.422772237042347   0.6794760987314773   0.3695407843355919   0.7549497990364407   0.8306013200848679   0.6272863969698881   0.579909633121213   0.736244269991129   0.7627571812455209   0.295185469203591   0.48491258375517926   0.7344386452278728   0.937164873863631   0.014003858220820306   0.5498834268881413   0.2168359538334019   0.41088061681246235   0.09623880895200809   0.00926805330261618   0.29228089929280693   0.6250404065431178   0.8062134323954078   0.027107946142560603   0.042467180471727574   0.20226816950077078   0.1267373336639305   0.6575671618069687   0.2875173814352869   0.37166684941590294   0.49945093669404245   0.07765752868575569   0.5512731114441578   0.608909668170382   0.20426546749045146   0.5927449449305765   0.816834466216285   0.6717447943067509   0.19026160926963115   0.04286151804243514   0.599998512382883   0.2608641774942886
0.09402280031762306   0.03359346473981896   0.3077176130900761   0.6358237709511708   0.28780936792221534   0.006485518597258354   0.2652504326183485   0.43355560145040006   0.1610720342582848   0.34891835679028965   0.9777330511830616   0.061888752034497105   0.6616210975642424   0.271260828104534   0.4264599397389038   0.4529790838641151   0.4573556300737909   0.6785158831739575   0.6096254735226189   0.7812342895573642   0.2670940208041597   0.6356543651315224   0.009626961139735818   0.5203701120630756   0.1730712204865367   0.6020609003917035   0.7019093480496598   0.8845463411119048   0.8852618525643213   0.595575381794445   0.4366589154313112   0.4509907396615047   0.7241898183060366   0.2466570250041554   0.45892586424824955   0.3891019876270076   0.0625687207417942   0.9753961968996214   0.03246592450934574   0.9361229037628924   0.6052130906680033   0.29688031372566387   0.4228404509867269   0.1548886142055283   0.33811906986384355   0.6612259485941415   0.4132134898469911   0.6345185021424528   0.16504784937730688   0.059165048202438064   0.7113041417973314   0.749972161030548   0.2797859968129855   0.463589666407993   0.2746452263660202   0.29898142136904327   0.555596178506949   0.21693264140383758   0.8157193621177706   0.9098794337420357   0.4930274577651547   0.24153644450421616   0.7832534376084249   0.9737565299791432
0.8878143670971514   0.9446561307785523   0.360412986621698   0.818867915773615   0.5496952972333079   0.2834301821844108   0.9471994967747069   0.1843494136311622   0.38464744785600097   0.2242651339819727   0.2358953549773756   0.4343772526006142   0.10486145104301549   0.7606754675739797   0.9612501286113554   0.13539583123157092   0.5492652725360665   0.5437428261701421   0.14553076649358482   0.22551639748953523   0.05623781477091182   0.30220638166592595   0.36227732888515995   0.25175986751039203   0.16842344767376038   0.3575502508873737   0.0018643422634619306   0.43289195173677714   0.6187281504404525   0.07412006870296291   0.05466484548875499   0.24854253810561494   0.23408070258445154   0.8498549347209902   0.8187694905113794   0.8141652855050008   0.12921925154143604   0.08917946714701047   0.857519361900024   0.6787694542734298   0.5799539790053695   0.5454366409768683   0.7119885954064392   0.4532530567838946   0.5237161642344577   0.24323025931094236   0.34971126652127926   0.20149318927350257   0.3552927165606973   0.8856800084235686   0.3478469242578173   0.7686012375367255   0.7365645661202448   0.8115599397206058   0.2931820787690623   0.5200586994311105   0.5024838635357932   0.9617050049996155   0.4744125882576829   0.7058934139261098   0.3732646119943572   0.8725255378526051   0.616893226357659   0.027123959652679958
0.7933106329889876   0.3270888968757368   0.9049046309512198   0.5738709028687854   0.26959446875452997   0.0838586375647944   0.5551933644299405   0.3723777135952828   0.9143017521938327   0.19817862914122575   0.20734644017212323   0.6037764760585573   0.17773718607358793   0.38661868942062   0.9141643614030609   0.08371777662744685   0.6752533225377947   0.42491368442100447   0.439751773145378   0.37782436270133707   0.30198871054343757   0.5523881465683994   0.8228585467877191   0.35070040304865713   0.5086780775544498   0.2252992496926626   0.9179539158364993   0.7768295001798717   0.23908360879991986   0.14144061212786818   0.3627605514065588   0.4044517865845889   0.32478185660608716   0.9432619829866424   0.15541411123443552   0.8006753105260316   0.1470446705324992   0.5566432935660224   0.24124974983137462   0.7169575338985847   0.4717913479947045   0.131729609145018   0.8014979766859966   0.3391331711972476   0.16980263745126695   0.5793414625766187   0.9786394298982776   0.9884327681485905   0.6611245598968171   0.35404221288395604   0.06068551406177833   0.21160326796871876   0.4220409510968972   0.21260160075608786   0.6979249626552195   0.8071514813841298   0.09725909449081006   0.2693396177694454   0.542510851420784   0.006476170858098262   0.9502144239583108   0.712696324203423   0.3012611015894094   0.2895186369595136
0.47842307596360634   0.580966715058405   0.49976312490341274   0.9503854657622659   0.3086204385123394   0.001625252481786382   0.5211236950051351   0.9619526976136754   0.6474958786155223   0.6475830395978304   0.4604381809433568   0.7503494296449567   0.22545492751862511   0.43498143884174245   0.7625132182881372   0.9431979482608268   0.12819583302781504   0.16564182107229705   0.2200023668673532   0.9367217774027286   0.1779814090695042   0.45294549686887403   0.9187412652779438   0.647203140443215   0.6995583331058979   0.8719787818104691   0.418978140374531   0.6968176746809491   0.39093789459355843   0.8703535293286826   0.8978544453693958   0.7348649770672737   0.7434420159780362   0.2227704897308523   0.4374162644260391   0.9845155474223171   0.517987088459411   0.7877890508891098   0.6749030461379019   0.0413175991614902   0.389791255431596   0.6221472298168128   0.4549006792705486   0.10459582175876164   0.21180984636209177   0.16920173294793875   0.5361594139926048   0.45739268131554667   0.5122515132561939   0.2972229511374697   0.11718127361807378   0.7605750066345975   0.12131361866263549   0.42686942180878706   0.21932682824867789   0.025710029567323885   0.37787160268459935   0.20409893207793475   0.7819105638226388   0.041194482145006865   0.8598845142251884   0.41630988118882495   0.107007517684737   0.9998768829835166
0.47009325879359243   0.7941626513720121   0.6521068384141884   0.895281061224755   0.25828341243150066   0.6249609184240734   0.11594742442158357   0.43788837990920837   0.7460318991753068   0.3277379672866037   0.9987661508035098   0.6773133732746108   0.6247182805126712   0.9008685454778166   0.779439322554832   0.6516033437072869   0.24684667782807188   0.6967696133998819   0.997528758732193   0.61040886156228   0.3869621636028835   0.28045973221105697   0.8905212410474561   0.6105319785787634   0.9168689048092911   0.4862970808390448   0.23841440263326769   0.7152509173540084   0.6585854923777904   0.8613361624149715   0.12246697821168412   0.2773625374448   0.9125535932024837   0.5335981951283677   0.12370082740817433   0.6000491641701892   0.2878353126898125   0.6327296496505511   0.34426150485334245   0.9484458204629023   0.040988634861740605   0.9359600362506693   0.34673274612114935   0.3380369589006222   0.6540264712588572   0.6555003040396122   0.4562115050736933   0.7275049803218587   0.737157566449566   0.16920322320056744   0.21779710244042558   0.012254062967850391   0.07857207407177556   0.307867060785596   0.09533012422874147   0.7348915255230504   0.16601848086929186   0.7742688656572283   0.9716292968205672   0.13484236135286118   0.8781831681794794   0.14153921600667718   0.6273677919672247   0.1863965408899589
0.8371945333177387   0.20557917975600798   0.2806350458460754   0.8483595819893367   0.18316806205888167   0.5500788757163957   0.8244235407723821   0.12085460166747795   0.44601049560931566   0.3808756525158283   0.6066264383319565   0.10860053869962756   0.3674384215375401   0.07300859173023228   0.5112963141032151   0.3737090131765772   0.20141994066824825   0.298739726073004   0.5396670172826479   0.238866651823716   0.32323677248876886   0.1572005100663268   0.9122992253154232   0.05247011093375707   0.4860422391710301   0.9516213303103188   0.6316641794693478   0.20411052894442033   0.3028741771121485   0.40154245459392307   0.8072406386969657   0.08325592727694239   0.8568636815028328   0.020666802078094793   0.20061420036500915   0.9746553885773148   0.4894252599652927   0.9476582103478625   0.6893178862617941   0.6009463754007377   0.2880053192970444   0.6489184842748585   0.1496508689791462   0.3620797235770217   0.9647685468082756   0.49171797420853175   0.23735164366372302   0.3096096126432646   0.47872630763724544   0.5400966438982129   0.6056874641943752   0.10549908369884425   0.17585213052509702   0.13855418930428984   0.7984468254974095   0.022243156421901857   0.3189884490222642   0.11788738722619505   0.5978326251324004   0.04758776784458702   0.8295631890569715   0.17022917687833253   0.9085147388706063   0.44664139244384937
0.541557869759927   0.521310692603474   0.75886386989146   0.08456166886682771   0.5767893229516515   0.029592718394942274   0.5215122262277371   0.7749520562235631   0.09806301531440602   0.4894960744967294   0.9158247620333618   0.6694529725247189   0.922210884789309   0.3509418851924395   0.11737793653595227   0.647209816102817   0.6032224357670448   0.23305449796624447   0.5195453114035519   0.59962204825823   0.7736592467100734   0.06282532108791195   0.6110305725329456   0.15298065581438064   0.23210137695014627   0.541514628484438   0.8521667026414855   0.06841898694755293   0.6553120539984948   0.5119219100894956   0.33065447641374845   0.2934669307239898   0.5572490386840887   0.022425835592766306   0.4148297143803866   0.624013958199271   0.6350381538947797   0.6714839504003268   0.29745177784443433   0.9768041420964539   0.03181571812773492   0.4384294524340823   0.7779064664408825   0.37718209383822393   0.2581564714176616   0.3756041313461704   0.1668758939079369   0.2242014380238433   0.026055094467515347   0.8340895028617324   0.31470919126645136   0.15578245107629038   0.37074304046902057   0.3221675927722368   0.9840547148527029   0.8623155203523005   0.8134940017849318   0.29974175717947044   0.5692250004723163   0.23830156215302964   0.17845584789015206   0.6282578067791437   0.27177322262788195   0.2614974200565757
0.14664012976241717   0.18982835434506135   0.4938667561869995   0.8843153262183518   0.8884836583447555   0.814224222998891   0.3269908622790626   0.6601138881945086   0.8624285638772402   0.9801347201371585   0.012281671012611203   0.5043314371182182   0.49168552340821964   0.6579671273649218   0.028226956159908265   0.6420159167659176   0.6781915216232878   0.35822537018545136   0.45900195568759194   0.40371435461288796   0.49973567373313577   0.7299675634063076   0.18722873305971   0.1422169345563122   0.3530955439707186   0.5401392090612464   0.6933619768727105   0.2579016083379604   0.46461188562596306   0.7259149860623553   0.3663711145936479   0.5977877201434518   0.6021833217487228   0.7457802659251968   0.3540894435810367   0.09345628302523373   0.11049779834050322   0.08781313856027495   0.32586248742112844   0.45144036625931616   0.4323062767172154   0.7295877683748236   0.8668605317335365   0.047726011646428215   0.9325706029840797   0.9996202049685159   0.6796317986738265   0.905509077090116   0.579475059013361   0.45948099590726965   0.986269821801116   0.6476074687521556   0.11486317338739799   0.7335660098449143   0.6198987072074681   0.04981974860870375   0.5126798516386751   0.9877857439197175   0.26580926362643137   0.9563634655834701   0.4021820532981719   0.8999726053594426   0.939946776205303   0.5049230993241539
0.9698757765809565   0.17038483698461898   0.07308624447176644   0.45719708767772566   0.037305173596876885   0.17076463201610304   0.3934544457979399   0.5516880105876096   0.45783011458351586   0.7112836361088334   0.4071846239968239   0.904080541835454   0.34296694119611787   0.9777176262639191   0.7872859167893558   0.8542607932267503   0.8302870895574427   0.9899318823442016   0.5214766531629245   0.8978973276432802   0.42810503625927077   0.08995927698475896   0.5815298769576215   0.3929742283191264   0.45822925967831424   0.91957444000014   0.5084436324858551   0.9357771406414007   0.4209240860814374   0.748809807984037   0.11498918668791515   0.3840891300537911   0.9630939714979215   0.03752617187520351   0.7078045626910913   0.4800085882183371   0.6201270303018037   0.0598085456112844   0.9205186459017354   0.6257477949915868   0.789839940744361   0.06987666326708285   0.39904199273881097   0.7278504673483066   0.3617349044850902   0.9799173862823239   0.8175121157811894   0.3348762390291802   0.903505644806776   0.060342946282183924   0.3090684832953344   0.39909909838777946   0.4825815587253386   0.311533138298147   0.19407929660741924   0.0150099683339884   0.5194875872274171   0.2740069664229435   0.48627473391632803   0.5350013801156513   0.8993605569256133   0.21419842081165907   0.5657560880145927   0.9092535851240645
0.10952061618125238   0.14432175754457624   0.16671409527578165   0.181403117775758   0.7477857116961621   0.16440437126225232   0.3492019794945922   0.8465268787465778   0.8442800668893863   0.10406142498006841   0.040133496199257816   0.4474277803587983   0.36169850816404764   0.7925282866819214   0.8460541995918386   0.4324178120248099   0.8422109209366306   0.5185213202589779   0.35977946567551056   0.8974164319091585   0.9428503640110173   0.30432289944731883   0.794023377660918   0.988162846785094   0.8333297478297649   0.16000114190274262   0.6273092823851364   0.806759729009336   0.08554403613360269   0.9955967706404902   0.27810730289054414   0.9602328502627583   0.24126396924421645   0.8915353456604219   0.23797380669128634   0.5128050699039599   0.8795654610801688   0.09900705897850046   0.39191960709944773   0.08038725787915003   0.03735454014353819   0.5804857387195226   0.032140141423937174   0.18297082596999145   0.09450417613252093   0.2761628392722037   0.23811676376301918   0.19480797918489742   0.26117442830275606   0.11616169736946107   0.6108074813778829   0.3880482501755614   0.17563039216915335   0.12056492672897079   0.3327001784873387   0.4278153999128031   0.9343664229249369   0.22902958106854893   0.09472637179605235   0.9150103300088431   0.054800961844768105   0.13002252209004844   0.7028067646966046   0.8346230721296931
0.017446421701229915   0.5495367833705259   0.6706666232726675   0.6516522461597016   0.922942245568709   0.2733739440983222   0.43254985950964825   0.45684426697480424   0.6617678172659529   0.15721224672886117   0.8217423781317654   0.06879601679924287   0.4861374250967996   0.036647319999890376   0.4890421996444267   0.6409806168864398   0.5517710021718627   0.8076177389313415   0.3943158278483743   0.7259702868775966   0.4969700403270946   0.677595216841293   0.6915090631517697   0.8913472147479035   0.4795236186258646   0.1280584334707671   0.020842439879102326   0.23969496858820183   0.5565813730571556   0.8546844893724449   0.5882925803694541   0.7828507016133975   0.8948135557912027   0.6974722426435837   0.7665502022376887   0.7140546848141547   0.4086761306944032   0.6608249226436933   0.27750800259326197   0.07307406792771494   0.8569051285225405   0.8532071837123518   0.8831921747448876   0.3471037810501183   0.35993508819544595   0.17561196687105884   0.19168311159311788   0.45575656630221484   0.8804114695695813   0.047553533400291746   0.17084067171401557   0.216061597714013   0.32383009651242567   0.19286904402784688   0.5825480913445614   0.4332108961006154   0.4290165407212229   0.49539680138426323   0.8159978891068728   0.7191562112864607   0.020340410026819765   0.8345718787405699   0.5384898865136108   0.6460821433587458
0.16343528150427925   0.9813646950282181   0.6552977117687232   0.29897836230862745   0.8035001933088333   0.8057527281571593   0.46361460017560524   0.8432217960064127   0.923088723739252   0.7581991947568675   0.2927739284615897   0.6271601982923997   0.5992586272268263   0.5653301507290206   0.7102258371170282   0.1939493021917842   0.17024208650560338   0.06993334934475737   0.8942279480101555   0.47479309090532346   0.1499016764787836   0.23536147060418747   0.35573806149654463   0.8287109475465777   0.9864663949745044   0.2539967755759694   0.7004403497278215   0.5297325852379502   0.18296620166567107   0.4482440474188102   0.23682574955221622   0.6865107892315376   0.2598774779264191   0.6900448526619427   0.9440518210906266   0.05935059093913797   0.6606188506995928   0.12471470193292218   0.2338259839735983   0.8654012887473538   0.4903767641939894   0.054781352588164814   0.33959803596344285   0.3906081978420303   0.3404750877152058   0.8194198819839773   0.9838599744668982   0.5618972502954527   0.35400869274070146   0.565423106408008   0.2834196247390767   0.03216466505750247   0.1710424910750304   0.11717905898919773   0.04659387518686047   0.3456538758259649   0.9111650131486113   0.42713420632725496   0.10254205409623394   0.28630328488682694   0.2505461624490185   0.3024195043943328   0.8687160701226356   0.42090199613947316
0.760169398255029   0.247638151806168   0.5291180341591928   0.03029379829744279   0.4196943105398233   0.42821826982219063   0.5452580596922946   0.4683965480019901   0.06568561779912185   0.8627951634141827   0.2618384349532179   0.4362318829444876   0.8946431267240915   0.7456161044249849   0.21524455976635745   0.09057800711852275   0.9834781135754802   0.31848189809773003   0.11270250567012349   0.8042747222316958   0.7329319511264617   0.01606239370339721   0.24398643554748783   0.38337272609222267   0.9727625528714325   0.7684242418972292   0.714868401388295   0.3530789277947799   0.5530682423316092   0.3402059720750386   0.16961034169600042   0.8846823797927897   0.48738262453248743   0.4774108086608559   0.9077719067427825   0.4484504968483022   0.592739497808396   0.7317947042358709   0.692527346976425   0.3578724897297794   0.6092613842329158   0.41331280613814086   0.5798248413063015   0.5535977674980835   0.8763294331064542   0.3972504124347437   0.3358384057588137   0.1702250414058609   0.9035668802350215   0.6288261705375144   0.6209700043705186   0.817146113611081   0.3504986379034123   0.28862019846247583   0.45135966267451827   0.9324637338182912   0.8631160133709249   0.8112093898016199   0.5435877559317358   0.48401323696998905   0.27037651556252895   0.07941468556574909   0.8510604089553108   0.1261407472402096
0.6611151313296132   0.6661018794276082   0.2712355676490092   0.572542979742126   0.7847856982231591   0.26885146699286455   0.9353971618901955   0.40231793833626517   0.8812188179881375   0.6400252964553501   0.3144271575196768   0.5851718247251841   0.5307201800847252   0.3514050979928742   0.8630674948451585   0.652708090906893   0.6676041667138003   0.5401957081912543   0.31947973891342274   0.16869485393690398   0.39722765115127134   0.4607810226255052   0.46841932995811203   0.04255410669669436   0.7361125198216582   0.794679143197897   0.19718376230910284   0.4700111269545683   0.951326821598499   0.5258276762050325   0.2617866004189074   0.06769318861830319   0.07010800361036154   0.8858023797496823   0.9473594428992306   0.482521363893119   0.5393878235256363   0.5343972817568081   0.08429194805407204   0.829813272986226   0.871783656811836   0.9942015735655538   0.7648122091406493   0.661118419049322   0.47455600566056466   0.5334205509400486   0.29639287918253726   0.6185643123526277   0.7384434858389065   0.7387414077421517   0.09920911687343444   0.14855318539805934   0.7871166642404075   0.21291373153711923   0.837422516454527   0.08085999677975615   0.717008660630046   0.32711135178743694   0.8900630735552965   0.5983386328866371   0.17762083710440962   0.7927140700306289   0.8057711255012244   0.7685253599004112
0.3058371802925736   0.798512496465075   0.040958916360575144   0.1074069408510891   0.8312811746320089   0.26509194552502646   0.7445660371780378   0.48884262849846144   0.0928376887931024   0.5263505377828748   0.6453569203046035   0.3402894431004021   0.3057210245526949   0.31343680624575554   0.8079344038500763   0.25942944632064596   0.588712363922649   0.9863254544583187   0.9178713302947799   0.6610908134340088   0.41109152681823935   0.19361138442768977   0.11210020479355541   0.8925654535335977   0.10525434652566576   0.39509888796261466   0.07114128843298026   0.7851585126825086   0.27397317189365683   0.13000694243758823   0.3265752512549424   0.29631588418404714   0.18113548310055444   0.6036564046547135   0.681218330950339   0.9560264410836451   0.8754144585478595   0.2902195984089579   0.8732839271002626   0.6965969947629991   0.2867020946252105   0.3038941439506393   0.9554125968054827   0.0355061813289903   0.8756105678069711   0.11028275952294951   0.8433123920119273   0.1429407277953926   0.7703562212813054   0.7151838715603348   0.772171103578947   0.357782215112884   0.49638304938764855   0.5851769291227465   0.44559585232400467   0.06146633092883685   0.31524756628709416   0.9815205244680332   0.7643775213736657   0.10543988984519179   0.4398331077392346   0.6913009260590752   0.8910935942734031   0.4088428950821927
0.1531310131140241   0.387406782108436   0.9356809974679203   0.3733367137532024   0.27752044530705294   0.27712402258548646   0.092368605455993   0.23039598595780977   0.5071642240257476   0.5619401510251516   0.32019750187704593   0.8726137708449258   0.010781174638098984   0.976763221902405   0.8746016495530412   0.811147439916089   0.6955336083510049   0.9952426974343719   0.11022412817937553   0.7057075500708971   0.2557005006117702   0.30394177137529665   0.21913053390597245   0.29686465498870446   0.10256948749774611   0.9165349892668607   0.2834495364380521   0.9235279412355021   0.8250490421906932   0.6394109666813742   0.1910809309820591   0.6931319552776923   0.31788481816494557   0.07747081565622262   0.8708834291050132   0.8205181844327666   0.3071036435268466   0.10070759375381758   0.996281779551972   0.009370744516677649   0.6115700351758417   0.10546489631944568   0.8860576513725964   0.30366319444578055   0.35586953456407155   0.801523124944149   0.6669271174666239   0.0067985394570760724   0.2533000470663255   0.8849881356772883   0.3834775810285718   0.083270598221574   0.4282510048756323   0.24557716899591409   0.19239665004651274   0.3901386429438817   0.11036618671068671   0.16810635333969148   0.32151322094149953   0.5696204585111151   0.80326254318384   0.0673987595858739   0.32523144138952764   0.5602497139944375
0.19169250800799834   0.9619338632664283   0.43917379001693124   0.25658651954865697   0.8358229734439268   0.1604107383222792   0.7722466725503073   0.24978798009158087   0.5825229263776013   0.27542260264499085   0.38876909152173544   0.1665173818700069   0.15427192150196903   0.02984543364907679   0.19637244147522268   0.7763787389261252   0.04390573479128232   0.8617390803093853   0.8748592205337231   0.20675828041501007   0.24064319160744224   0.7943403207235115   0.5496277791441955   0.6465085664205726   0.048950683599443906   0.8324064574570832   0.11045398912726427   0.3899220468719156   0.21312771015551712   0.671995719134804   0.338207316576957   0.14013406678033474   0.6306047837779158   0.39657311648981314   0.9494382250552216   0.9736166849103278   0.4763328622759468   0.3667276828407363   0.7530657835799989   0.19723794598420266   0.4324271274846645   0.504988602531351   0.8782065630462758   0.9904796655691925   0.19178393587722223   0.7106482818078396   0.32857878390208023   0.34397109914862   0.14283325227777832   0.8782418243507564   0.21812479477481597   0.9540490522767043   0.9297055421222612   0.2062461052159524   0.8799174781978589   0.8139149854963696   0.2991007583443454   0.8096729887261392   0.9304792531426374   0.8402983005860417   0.8227678960683986   0.44294530588540293   0.17741346956263854   0.6430603546018391
0.3903407685837341   0.9379567033540519   0.2992069065163628   0.6525806890326464   0.1985568327065119   0.22730842154621234   0.9706281226142826   0.3086095898840265   0.05572358042873355   0.3490665971954559   0.7525033278394665   0.35456053760732215   0.12601803830647235   0.14282049197950353   0.8725858496416076   0.5406455521109526   0.8269172799621269   0.33314750325336423   0.9421065964989702   0.7003472515249107   0.004149383893728371   0.8902021973679614   0.7646931269363316   0.05728689692307171   0.6138086153099942   0.9522454940139093   0.46548622041996884   0.4047062078904252   0.41525178260348233   0.724937072467697   0.49485809780568635   0.09609661800639875   0.3595282021747488   0.3758704752722411   0.7423547699662199   0.7415360803990766   0.23351016386827644   0.23304998329273757   0.8697689203246122   0.2008905282881241   0.4065928839061495   0.8999024800393733   0.9276623238256421   0.5005432767632133   0.40244350001242113   0.009700282671412019   0.1629691968893104   0.4432563798401416   0.7886348847024268   0.05745478865750265   0.6974829764693415   0.038550171949716376   0.3733831020989445   0.33251771618980563   0.2026248786636552   0.9424535539433176   0.013854899924195703   0.9566472409175645   0.4602701086974354   0.200917473544241   0.7803447360559193   0.723597257624827   0.5905011883728232   0.00002694525611691024
0.37375185214976975   0.8236947775854536   0.6628388645471811   0.4994836684929036   0.9713083521373487   0.8139944949140416   0.4998696676578707   0.05622728865276199   0.18267346743492177   0.756539706256539   0.8023866911885291   0.01767711670304561   0.8092903653359773   0.42402199006673336   0.5997618125248739   0.07522356275972798   0.7954354654117816   0.4673747491491688   0.13949170382743856   0.874306089215487   0.015090729355862309   0.7437774915243419   0.5489905154546154   0.87427914395937   0.6413388772060925   0.9200827139388883   0.8861516509074343   0.37479547546646647   0.6700305250687439   0.10608821902484666   0.38628198324956353   0.31856818681370447   0.48735705763382214   0.34954851276830773   0.5838952920610344   0.30089107011065885   0.6780666922978449   0.9255265227015744   0.9841334795361604   0.22566750735093088   0.8826312268860633   0.45815177355240555   0.8446417757087219   0.3513614181354439   0.867540497530201   0.7143742820280636   0.2956512602541065   0.47708227417607385   0.22620162032410845   0.7942915680891754   0.4094996093466722   0.10228679870960738   0.5561710952553646   0.6882033490643288   0.023217626097108642   0.7837186118959029   0.06881403762154242   0.338654836296021   0.43932233403607424   0.48282754178524406   0.39074734532369754   0.41312831359444663   0.45518885449991386   0.2571600344343132
0.5081161184376343   0.954976540042041   0.610547078791192   0.9057986162988693   0.6405756209074333   0.24060225801397742   0.31489581853708554   0.4287163421227954   0.4143740005833248   0.446310689924802   0.9053962091904133   0.32642954341318803   0.8582029053279603   0.7581073408604733   0.8821785830933047   0.5427109315172851   0.7893888677064178   0.41945250456445227   0.4428562490572304   0.059883389732041055   0.39864152238272027   0.006324190970005638   0.9876673945573166   0.8027233552977279   0.8905254039450861   0.05134765092796456   0.3771203157661246   0.8969247389988586   0.24994978303765278   0.8107453929139872   0.06222449722903906   0.46820839687606325   0.835575782454328   0.3644347029891852   0.15682828803862572   0.14177885346287525   0.9773728771263677   0.6063273621287119   0.27464970494532104   0.5990679219455901   0.18798400941994986   0.18687485756425962   0.8317934558880906   0.5391845322135491   0.7893424870372295   0.18055066659425398   0.844126061330774   0.7364611769158212   0.8988170830921435   0.12920301566628942   0.4670057455646494   0.8395364379169625   0.6488673000544908   0.31845762275230227   0.40478124833561036   0.3713280410408993   0.8132915176001627   0.9540229197631171   0.2479529602969846   0.22954918757802406   0.835918640473795   0.34769555763440524   0.9733032553516636   0.6304812656324339
0.6479346310538452   0.16082070007014562   0.141509799463573   0.09129673341888478   0.8585921440166157   0.9802700334758916   0.297383738132799   0.35483555650306353   0.9597750609244721   0.8510670178096023   0.8303779925681496   0.515299118586101   0.31090776086998134   0.5326093950573   0.42559674423253924   0.1439710775452017   0.4976162432698186   0.578586475294183   0.17764378393555463   0.9144218899671777   0.6616976027960235   0.23089091765977768   0.20434052858389107   0.28394062433474376   0.013762971742178371   0.07007021758963206   0.06283072912031806   0.19264389091585898   0.15517082772556276   0.08980018411374041   0.7654469909875191   0.8378083344127955   0.19539576680109064   0.23873316630413818   0.9350689984193694   0.32250921582669445   0.8844880059311093   0.7061237712468382   0.5094722541868302   0.17853813828149276   0.38687176266129064   0.1275372959526553   0.33182847025127554   0.2641162483143151   0.7251741598652671   0.8966463782928776   0.1274879416673845   0.9801756239795714   0.7114111881230888   0.8265761607032456   0.06465721254706644   0.7875317330637124   0.556240360397526   0.7367759765895051   0.2992102215595474   0.9497233986509169   0.36084459359643534   0.49804281028536695   0.36414122314017794   0.6272141828242226   0.47635658766532607   0.7919190390385288   0.8546689689533478   0.4486760445427298
0.0894848250040354   0.6643817430858735   0.5228404987020722   0.18455979622841467   0.3643106651387683   0.7677353647929959   0.39535255703468763   0.2043841722488433   0.6528994770156795   0.9411592040897503   0.3306953444876212   0.41685243918513093   0.09665911661815357   0.20438322750024512   0.03148512292807384   0.46712904053421395   0.7358145230217182   0.7063404172148782   0.6673438997878959   0.8399148577099914   0.25945793535639217   0.9144213781763494   0.8126749308345482   0.3912388131672616   0.16997311035235677   0.2500396350904759   0.28983443213247606   0.20667901693884694   0.8056624452135884   0.4823042702974801   0.8944818750977884   0.0022948446900036305   0.1527629681979089   0.5411450662077297   0.5637865306101671   0.5854424055048727   0.05610385157975535   0.33676183870748466   0.5323014076820933   0.1183133649706588   0.3202893285580371   0.6304214214926065   0.8649575078941975   0.2783985072606674   0.060831393201644955   0.7160000433162571   0.05228257705964921   0.8871596940934058   0.8908582828492881   0.4659604082257812   0.7624481449271732   0.6804806771545588   0.08519583763569971   0.9836561379283012   0.8679662698293847   0.6781858324645552   0.9324328694377908   0.44251107172057136   0.30417973921921765   0.0927434269596825   0.8763290178580354   0.10574923301308671   0.7718783315371243   0.9744300619890237
0.5560396892999984   0.4753278115204802   0.9069208236429269   0.6960315547283563   0.4952082960983534   0.7593277682042231   0.8546382465832777   0.8088718606349505   0.6043500132490652   0.2933673599784419   0.0921901016561045   0.12839118348039166   0.5191541756133655   0.30971122205014073   0.2242238318267197   0.4502053510158364   0.5867213061755747   0.8672001503295693   0.9200440926075021   0.3574619240561539   0.7103922883175392   0.7614509173164826   0.14816576107037777   0.3830318620671302   0.15435259901754092   0.2861231057960024   0.2412449374274509   0.6870003073387739   0.6591443029191876   0.5267953375917793   0.3866066908441732   0.8781284467038234   0.05479428967012235   0.23342797761333747   0.29441658918806873   0.7497372632234317   0.5356401140567569   0.9237167555631968   0.07019275736134903   0.2995319122075953   0.9489188078811822   0.056516605233627386   0.15014866475384694   0.9420699881514414   0.23852651956364296   0.29506568791714477   0.001982903683469179   0.5590381260843111   0.08417392054610205   0.008942582121142314   0.7607379662560183   0.8720378187455373   0.4250296176269145   0.482147244529363   0.37413127541184504   0.9939093720417139   0.37023532795679215   0.2487192669160255   0.07971468622377634   0.24417210881828222   0.8345952139000353   0.32500251135282876   0.009521928862427309   0.944640196610687
0.8856764060188531   0.26848590611920137   0.8593732641085804   0.002570208459245619   0.6471498864552101   0.9734202182020566   0.8573903604251112   0.44353208237493447   0.562975965909108   0.9644776360809143   0.09665239416909288   0.5714942636293971   0.13794634828219354   0.48233039155155133   0.7225211187572478   0.5775848915876832   0.7677110203254014   0.23361112463552583   0.6428064325334715   0.33341278276940106   0.9331158064253661   0.908608613282697   0.6332845036710442   0.3887725861587141   0.04743940040651302   0.6401227071634957   0.7739112395624638   0.38620237769946847   0.4002895139513029   0.666702488961439   0.9165208791373527   0.942670295324534   0.8373135480421948   0.7022248528805247   0.8198684849682598   0.3711760316951368   0.6993671997600013   0.2198944613289734   0.09734736621101193   0.7935911401074536   0.9316561794345999   0.9862833366934476   0.45454093367754045   0.46017835733805246   0.9985403730092338   0.07767472341075048   0.8212564300064963   0.0714057711793384   0.9511009726027208   0.4375520162472548   0.047345190444032445   0.6852033934798699   0.5508114586514179   0.7708495272858157   0.1308243113066798   0.742533098155336   0.7134979106092231   0.068624674405291   0.31095582633842006   0.37135706646019917   0.014130710849221772   0.8487302130763176   0.2136084601274081   0.5777659263527456
0.0824745314146219   0.8624468763828701   0.7590675264498676   0.11758756901469317   0.08393415840538813   0.7847721529721196   0.9378110964433714   0.04618179783535477   0.13283318580266737   0.3472201367248648   0.890465905999339   0.36097840435548484   0.5820217271512496   0.576370609439049   0.7596415946926591   0.6184453062001488   0.8685238165420265   0.5077459350337581   0.4486857683542391   0.2470882397399497   0.8543931056928047   0.6590157219574404   0.23507730822683098   0.669322313387204   0.7719185742781828   0.7965688455745704   0.47600978177696335   0.5517347443725109   0.6879844158727947   0.011796692602450793   0.5381986853335919   0.5055529465371561   0.5551512300701273   0.664576555877586   0.647732779334253   0.1445745421816713   0.9731295029188778   0.08820594643853695   0.8880911846415939   0.5261292359815224   0.1046056863768513   0.5804600114047789   0.4394054162873548   0.27904099624157275   0.2502125806840466   0.9214442894473385   0.2043281080605238   0.6097186828543687   0.4782940064058638   0.12487544387276807   0.7283183262835604   0.05798393848185781   0.7903095905330692   0.11307875127031727   0.1901196409499685   0.5524309919447017   0.2351583604629418   0.4485021953927313   0.5423868616157155   0.4078564497630304   0.262028857544064   0.3602962489541943   0.6542956769741216   0.881727213781508
0.15742317116721272   0.7798362375494154   0.2148902606867668   0.6026862175399352   0.9072105904831661   0.858391948102077   0.010562152626243016   0.9929675346855665   0.4289165840773023   0.7335165042293089   0.2822438263426826   0.9349835962037087   0.6386069935442332   0.6204377529589916   0.09212418539271407   0.382552604259007   0.4034486330812914   0.17193555756626036   0.5497373237769986   0.9746961544959766   0.14141977553722743   0.811639308612066   0.895441646802877   0.09296894071446865   0.9839966043700147   0.031803071062650595   0.6805513861161102   0.4902827231745334   0.0767860138868486   0.1734111229605736   0.6699892334898672   0.4973151884889669   0.6478694298095462   0.4398946187312647   0.38774540714718464   0.5623315922852582   0.009262436265313005   0.8194568657722731   0.29562122175447053   0.17977898802625114   0.6058138031840216   0.6475213082060127   0.7458838979774719   0.20508283353027454   0.4643940276467941   0.8358819995939466   0.8504422511745949   0.11211389281580587   0.4803974232767794   0.804078928531296   0.16989086505848472   0.6218311696412724   0.40361140938993084   0.6306678055707224   0.49990163156861755   0.12451598115230554   0.7557419795803846   0.19077318683945776   0.11215622442143292   0.5621843888670474   0.7464795433150716   0.3713163210671847   0.8165350026669623   0.3824054008407962
0.14066574013105002   0.723795012861172   0.07065110468949043   0.17732256731052168   0.6762717124842559   0.8879130132672254   0.2202088535148955   0.06520867449471582   0.19587428920747646   0.08383408473592935   0.05031798845641076   0.44337750485344335   0.7922628798175456   0.4531662791652069   0.5504163568877932   0.31886152370113785   0.03652090023716108   0.26239309232574914   0.4382601324663603   0.7566771348340905   0.2900413569220895   0.8910767712585644   0.6217251297993979   0.3742717339932943   0.1493756167910395   0.1672817583973924   0.5510740251099074   0.19694916668277257   0.4731039043067836   0.279368745130167   0.330865171595012   0.13174049218805678   0.27722961509930716   0.19553466039423767   0.2805471831386012   0.6883629873346134   0.4849667352817615   0.7423683812290307   0.730130826250808   0.3695014636334756   0.44844583504460045   0.4799752889032816   0.29187069378444774   0.6128243287993851   0.15840447812251093   0.5888985176447171   0.6701455639850498   0.23855259480609084   0.009028861331471419   0.4216167592473247   0.11907153887514232   0.04160342812331825   0.5359249570246878   0.1422480141171577   0.7882063672801303   0.9098629359352615   0.25869534192538063   0.9467133537229201   0.5076591841415291   0.2214999486006481   0.7737286066436191   0.2043449724938893   0.7775283578907211   0.8519984849671726
0.3252827715990187   0.7243696835906077   0.4856576641062733   0.23917415616778745   0.1668782934765078   0.13547116594589056   0.8155121001212235   0.0006215613616966076   0.15784943214503636   0.7138544066985658   0.6964405612460812   0.9590181332383784   0.6219244751203485   0.5716063925814081   0.9082341939659508   0.04915519730311687   0.3632291331949679   0.6248930388584881   0.4005750098244218   0.8276552487024688   0.5895005265513488   0.4205480663645988   0.6230466519337007   0.9756567637352963   0.2642177549523301   0.696178382773991   0.1373889878274274   0.7364826075675088   0.09733946147582231   0.5607072168281005   0.3218768877062039   0.7358610462058122   0.939490029330786   0.8468528101295346   0.6254363264601227   0.7768429129674339   0.31756555421043736   0.2752464175481265   0.7172021324941719   0.727687715664317   0.9543364210154694   0.6503533786896384   0.31662712266975007   0.9000324669618482   0.3648358944641207   0.22980531232503965   0.6935804707360493   0.9243757032265519   0.10061813951179056   0.5336269295510486   0.556191482908622   0.18789309565904314   0.0032786780359682563   0.9729197127229481   0.23431459520241807   0.45203204945323094   0.0637886487051823   0.12606690259341344   0.6088782687422953   0.675189136485797   0.7462230944947449   0.850820485045287   0.8916761362481235   0.94750142082148
0.7918866734792754   0.2004671063556485   0.5750490135783735   0.04746895385963189   0.4270507790151548   0.9706617940306088   0.881468542842324   0.12309325063307995   0.32643263950336426   0.43703486447956025   0.3252770599337021   0.9352001549740369   0.323153961467396   0.46411515175661217   0.09096246473128404   0.4831681055208059   0.2593653127622137   0.3380482491631987   0.4820841959889887   0.8079789690350089   0.5131422182674688   0.4872277641179118   0.5904080597408652   0.8604775482135287   0.7212555447881933   0.2867606577622633   0.015359046162491773   0.8130085943538968   0.29420476577303845   0.31609886373165447   0.13389050332016772   0.6899153437208169   0.9677721262696742   0.8790639992520942   0.8086134433864656   0.7547151887467801   0.6446181648022782   0.4149488474954821   0.7176509786551816   0.2715470832259742   0.38525285204006454   0.07690059833228338   0.23556678266619288   0.4635681141909654   0.8721106337725958   0.5896728342143716   0.6451587229253277   0.6030905659774366   0.15085508898440253   0.30291217645210833   0.6297996767628359   0.7900819716235398   0.856650323211364   0.9868133127204538   0.4959091734426682   0.10016662790272285   0.8888781969416898   0.10774931346835964   0.6872957300562026   0.34545143915594273   0.24426003213941158   0.6928004659728776   0.969644751401021   0.07390435592996855
0.8590071800993471   0.6158998676405941   0.7340779687348281   0.6103362417390032   0.9868965463267513   0.02622703342622256   0.08891924580950047   0.007245675761566581   0.8360414573423487   0.7233148569741142   0.45911956904666457   0.21716370413802683   0.9793911341309847   0.7365015442536603   0.9632103956039963   0.11699707623530398   0.09051293718929483   0.6287522307853007   0.27591466554779376   0.7715456370793612   0.8462529050498833   0.9359517648124231   0.30626991414677274   0.6976412811493927   0.9872457249505362   0.320051897171829   0.5721919454119446   0.08730503941038949   0.0003491786237849806   0.29382486374560646   0.4832726996024441   0.0800593636488229   0.16430772128143628   0.5705100067714922   0.024153130555779567   0.862895659510796   0.18491658715045162   0.8340084625178319   0.060942734951783206   0.7458985832754921   0.09440364996115679   0.2052562317325311   0.7850280694039894   0.9743529461961309   0.24815074491127356   0.2693044669201079   0.4787581552572167   0.27671166504673816   0.26090501996073734   0.9492525697482789   0.9065662098452721   0.1894066256363487   0.26055584133695237   0.6554277060026724   0.42329351024282796   0.10934726198752578   0.09624812005551608   0.08491769923118023   0.3991403796870484   0.2464516024767297   0.9113315329050644   0.25090923671334836   0.3381976447352652   0.5005530192012376
0.8169278829439077   0.045653004980817286   0.5531695753312758   0.5262000730051067   0.5687771380326341   0.7763485380607094   0.07441142007405907   0.24948840795836857   0.3078721180718968   0.8270959683124305   0.16784521022878698   0.060081782322019876   0.04731627673494443   0.17166826230975804   0.744551699985959   0.9507345203344941   0.9510681566794283   0.08675056307857781   0.3454113202989106   0.7042829178577644   0.03973662377436387   0.8358413263652295   0.007213675563645391   0.20372989865652677   0.22280874083045618   0.7901883213844122   0.45404410023236963   0.6775298256514201   0.654031602797822   0.013839783323702767   0.37963268015831053   0.42804141769305143   0.3461594847259253   0.1867438150112723   0.21178746992952358   0.3679596353710316   0.29884320799098085   0.01507555270151425   0.4672357699435646   0.4172251150365375   0.3477750513115525   0.9283249896229364   0.12182444964465397   0.7129421971787732   0.30803842753718863   0.092483663257707   0.11461077408100859   0.5092122985222464   0.08522968670673245   0.3022953418732949   0.660566673848639   0.8316824728708263   0.4311980839089104   0.2884555585495921   0.2809339936903284   0.4036410551777749   0.0850385991829851   0.1017117435383198   0.06914652376080484   0.03568141980674331   0.7861953911920042   0.08663619083680556   0.6019107538172402   0.6184563047702059
0.43842033988045176   0.15831120121386913   0.4800863041725863   0.9055141075914327   0.1303819123432631   0.06582753795616211   0.36547553009157774   0.3963018090691864   0.045152225636530645   0.7635321960828673   0.7049088562429388   0.56461933619836   0.6139541417276203   0.47507663753327517   0.42397486255261035   0.16097828102058515   0.5289155425446351   0.37336489399495537   0.3548283387918055   0.12529686121384181   0.7427201513526309   0.2867287031581498   0.7529175849745652   0.506840556443636   0.30429981147217916   0.12841750194428067   0.27283128080197894   0.6013264488522033   0.1739178991289161   0.06258996398811856   0.9073557507104012   0.20502463978301694   0.12876567349238546   0.2990577679052513   0.20244689446746247   0.6404053035846569   0.5148115317647652   0.8239811303719762   0.7784720319148521   0.47942702256407177   0.98589598922013   0.4506162363770208   0.4236436931230466   0.35413016135022996   0.2431758378674991   0.163887533218871   0.6707261081484814   0.847289604906594   0.93887602639532   0.035470031274590336   0.39789482734650244   0.24596315605439065   0.7649581272664039   0.9728800672864718   0.49053907663610125   0.040938516271373716   0.6361924537740183   0.6738222993812204   0.2880921821686388   0.4005332126867168   0.1213809220092532   0.8498411690092443   0.5096201502537867   0.921106190122645
0.13548493278912316   0.3992249326322235   0.08597645713074004   0.566976028772415   0.892309094921624   0.2353373994133525   0.41525034898225865   0.7196864238658212   0.9534330685263042   0.19986736813876216   0.017355521635756193   0.4737232678114305   0.1884749412599003   0.22698730085229038   0.526816444999655   0.43278475154005674   0.5522824874858819   0.55316500147107   0.23872426283101617   0.032251538853339964   0.4309015654766287   0.7033238324618256   0.7291041125772295   0.11114534873069494   0.29541663268750556   0.30409889982960214   0.6431276554464894   0.5441693199582799   0.4031075377658815   0.06876150041624965   0.22787730646423082   0.8244828960924587   0.4496744692395774   0.8688941322774875   0.2105217848284746   0.35075962828102825   0.26119952797967705   0.6419068314251971   0.6837053398288196   0.9179748767409714   0.7089170404937951   0.08874182995412717   0.4449810769978035   0.8857233378876315   0.27801547501716645   0.38541799749230155   0.715876964420574   0.7745779891569365   0.9825988423296609   0.08131909766269942   0.07274930897408452   0.2304086691986567   0.5794913045637794   0.012557597246449776   0.8448720025098537   0.405925773106198   0.129816835324202   0.1436634649689623   0.6343502176813791   0.05516614482516976   0.8686173073445249   0.5017566335437652   0.9506448778525595   0.1371912680841983
0.15970026685072974   0.413014803589638   0.5056638008547559   0.25146793019656677   0.8816847918335633   0.02759680609733646   0.7897868364341819   0.4768899410396302   0.8990859495039024   0.946277708434637   0.7170375274600974   0.24648127184097351   0.31959464494012313   0.9337201111881872   0.8721655249502437   0.8405554987347755   0.1897778096159211   0.790056646219225   0.2378153072688646   0.7853893539096057   0.3211605022713962   0.2883000126754598   0.28717042941630516   0.6481980858254075   0.16146023542066645   0.8752852090858217   0.7815066285615493   0.3967301556288407   0.2797754435871031   0.8476884029884854   0.9917197921273674   0.9198402145892105   0.3806894940832007   0.9014106945538483   0.2746822646672699   0.6733589427482369   0.06109484914307755   0.967690583365661   0.40251673971702623   0.8328034440134614   0.8713170395271564   0.17763393714643605   0.16470143244816163   0.047414090103855694   0.5501565372557602   0.8893339244709763   0.8775310030318564   0.3992160042784482   0.38869630183509374   0.014048715385154474   0.09602437447030716   0.0024858486496075454   0.10892085824799062   0.16636031239666915   0.10430458234293984   0.08264563406039709   0.72823136416479   0.26494961784282084   0.82962231767567   0.4092866913121601   0.6671365150217125   0.29725903447715984   0.4271055779586437   0.5764832472986987
0.795819475494556   0.1196250973307238   0.2624041455104821   0.5290691571948429   0.24566293823879579   0.23029117285974754   0.38487314247862564   0.12985315291639477   0.8569666364037021   0.21624245747459306   0.2888487680083185   0.12736730426678722   0.7480457781557114   0.04988214507792391   0.18454418566537864   0.044721670206390125   0.019814413990921428   0.7849325272351031   0.35492186798970876   0.63543497889423   0.35267789896920904   0.4876734927579432   0.927816290031065   0.05895173159553133   0.556858423474653   0.3680483954272194   0.665412144520583   0.5298825744006883   0.3111954852358572   0.13775722256747186   0.2805390020419573   0.4000294214842936   0.4542288488321552   0.9215147650928788   0.9916902340336389   0.2726621172175064   0.7061830706764438   0.8716326200149549   0.8071460483682602   0.22794044701111627   0.6863686566855224   0.08670009277985184   0.4522241803785515   0.5925054681168862   0.3336907577163134   0.5990266000219087   0.5244078903474865   0.533553736521355   0.7768323342416603   0.23097820459468923   0.8589957458269034   0.003671162120666576   0.4656368490058031   0.09322098202721738   0.5784567437849462   0.603641740636373   0.011408000173647915   0.17170621693433857   0.5867665097513073   0.3309796234188666   0.3052249294972041   0.3000735969193837   0.7796204613830471   0.10303917640775033
0.6188562728116818   0.21337350413953182   0.3273962810044956   0.5105337082908641   0.28516551509536836   0.6143469041176232   0.8029883906570091   0.9769799717695091   0.5083331808537079   0.38336869952293395   0.9439926448301057   0.9733088096488426   0.042696331847904855   0.2901477174957166   0.3655359010451596   0.3696670690124696   0.03128833167425694   0.11844150056137802   0.7787693912938524   0.038687445593603   0.7260634021770528   0.8183679036419943   0.9991489299108053   0.9356482691858526   0.10720712936537112   0.6049943995024625   0.6717526489063097   0.4251145608949886   0.8220416142700028   0.9906474953848393   0.8687642582493006   0.44813458912547943   0.3137084334162948   0.6072787958619054   0.9247716134191949   0.47482577947663684   0.27101210156838995   0.31713107836618876   0.5592357123740352   0.10515871046416726   0.239723769894133   0.19868957780481075   0.780466321080183   0.06647126487056426   0.5136603677170801   0.3803216741628164   0.7813173911693777   0.1308229956847116   0.40645323835170905   0.7753272746603539   0.10956474226306796   0.705708434789723   0.5844116240817063   0.7846797792755146   0.2408004840137674   0.2575738456642436   0.2707031906654115   0.17740098341360921   0.3160288705945726   0.7827480661876067   0.9996910890970215   0.8602699050474204   0.7567931582205373   0.6775893557234395
0.7599673192028885   0.6615803272426097   0.9763268371403544   0.6111180908528752   0.24630695148580836   0.2812586530797933   0.1950094459709767   0.4802950951681636   0.8398537131340993   0.5059313784194394   0.08544470370790873   0.7745866603784406   0.255442089052393   0.7212515991439248   0.8446442196941413   0.517012814714197   0.9847388983869816   0.5438506157303156   0.5286153490995688   0.7342647485265903   0.98504780928996   0.6835807106828952   0.7718221908790315   0.056675392803150856   0.2250804900870715   0.022000383440285463   0.7954953537386771   0.44555730195027565   0.9787735386012631   0.7407417303604922   0.6004859077677004   0.965262206782112   0.13891982546716383   0.23481035194105276   0.5150412040597917   0.19067554640367143   0.8834777364147708   0.5135587527971279   0.6703969843656504   0.6736627316894744   0.8987388380277892   0.9697081370668124   0.14178163526608162   0.939397983162884   0.9136910287378293   0.28612742638391714   0.36995944438705014   0.8827225903597332   0.6886105386507577   0.2641270429436317   0.574464090648373   0.43716528840945756   0.7098370000494946   0.5233853125831396   0.9739781828806726   0.4719030816273455   0.5709171745823307   0.28857496064208676   0.45893697882088086   0.2812275352236741   0.6874394381675599   0.7750162078449588   0.7885399944552305   0.6075648035341997
0.7887006001397707   0.8053080707781465   0.6467583591891488   0.6681668203713156   0.8750095714019415   0.5191806443942294   0.27679891480209873   0.7854442300115824   0.1863990327511838   0.25505360145059763   0.7023348241537257   0.34827894160212486   0.47656203270168923   0.7316682888674582   0.7283566412730531   0.8763758599747793   0.9056448581193585   0.44309332822537134   0.2694196624521722   0.5951483247511052   0.2182054199517985   0.6680771203804126   0.4808796679969417   0.9875835212169055   0.4295048198120278   0.862769049602266   0.8341213088077929   0.3194167008455899   0.5544952484100863   0.34358840520803663   0.5573223940056942   0.5339724708340075   0.3680962156589025   0.088534803757439   0.8549875698519684   0.1856935292318826   0.8915341829572133   0.3568665148899809   0.1266309285789154   0.3093176692571033   0.9858893248378549   0.9137731866646095   0.8572112661267433   0.7141693445059981   0.7676839048860563   0.245696066284197   0.3763315981298015   0.7265858232890926   0.3381790850740285   0.382927016681931   0.5422102893220087   0.40716912244350273   0.7836838366639421   0.03933861147389434   0.9848878953163145   0.8731966516094952   0.41558762100503965   0.9508038077164553   0.12990032546434602   0.6875031223776127   0.5240534380478264   0.5939372928264745   0.0032693968854306237   0.3781854531205094
0.5381641132099716   0.680164106161865   0.14605813075868743   0.6640161086145113   0.7704802083239153   0.43446803987766797   0.7697265326288859   0.9374302853254187   0.4323011232498868   0.051541023195736946   0.22751624330687728   0.530261162881916   0.6486172865859446   0.012202411721842606   0.24262834799056276   0.6570645112724207   0.23302966558090493   0.06139860400538726   0.11272802252621675   0.969561388894808   0.7089762275330785   0.4674613111789128   0.10945862564078612   0.5913759357742987   0.17081211432310697   0.7872972050170478   0.9634004948820987   0.9273598271597874   0.40033190599919166   0.3528291651393799   0.1936739622532128   0.9899295418343688   0.9680307827493049   0.30128814194364295   0.9661577189463355   0.4596683789524527   0.31941349616336023   0.28908573022180034   0.7235293709557727   0.802603867680032   0.08638383058245531   0.2276871262164131   0.610801348429556   0.8330424787852239   0.37740760304937676   0.7602258150375003   0.5013427227887699   0.2416665430109252   0.20659548872626982   0.9729286100204525   0.5379422279066711   0.3143067158511378   0.8062635827270781   0.6200994448810725   0.34426826565345836   0.324377174016769   0.8382327999777732   0.3188113029374296   0.37811054670712285   0.8647087950643163   0.518819303814413   0.02972557271562924   0.6545811757513501   0.06210492738428433
0.4324354732319577   0.8020384464992162   0.04377982732179413   0.22906244859906041   0.05502787018258094   0.04181263146171586   0.5424371045330243   0.9873959055881353   0.8484323814563112   0.06888402144126342   0.00449487662635309   0.6730891897369975   0.042168798729232994   0.4487845765601909   0.6602266109728947   0.3487120157202284   0.2039359987514597   0.1299732736227613   0.28211606426577185   0.4840032206559121   0.6851166949370467   0.10024770090713205   0.6275348885144217   0.42189829327162776   0.252681221705089   0.2982092544079159   0.5837550611926275   0.19283584467256734   0.19765335152250804   0.2563966229462   0.04131795665960329   0.20543993908443212   0.3492209700661969   0.18751260150493662   0.0368230800332502   0.5323507493474346   0.3070521713369639   0.7387280249447458   0.3765964690603555   0.18363873362720623   0.10311617258550418   0.6087547513219844   0.09448040479458368   0.6996355129712941   0.4179994776484575   0.5085070504148524   0.466945516280162   0.27773721969966636   0.16531825594336852   0.21029779600693652   0.8831904550875345   0.084901375027099   0.9676649044208605   0.9539011730607365   0.8418724984279311   0.8794614359426669   0.6184439343546636   0.7663885715557999   0.8050494183946809   0.3471106865952322   0.31139176301769966   0.02766054661105414   0.42845294933432543   0.16347195296802597
0.2082755904321955   0.4189057952890697   0.33397254453974173   0.46383643999673185   0.790276112783738   0.9103987448742172   0.8670270282595798   0.1860992202970655   0.6249578568403695   0.7001009488672807   0.9838365731720453   0.10119784526996649   0.657292952419509   0.7461997758065443   0.1419640747441142   0.22173640932729963   0.03884901806484542   0.9798112042507443   0.3369146563494333   0.8746257227320674   0.7274572550471458   0.9521506576396902   0.9084617070151079   0.7111537697640414   0.5191816646149502   0.5332448623506205   0.5744891624753661   0.24731732976730955   0.7289055518312122   0.6228461174764033   0.7074621342157863   0.061218109470244066   0.10394769499084273   0.9227451686091226   0.723625561043741   0.9600202642002775   0.4466547425713337   0.17654539280257833   0.5816614862996268   0.738283854872978   0.40780572450648833   0.19673418855183397   0.2447468299501935   0.8636581321409106   0.6803484694593426   0.24458353091214377   0.33628512293508567   0.15250436237686915   0.16116680484439233   0.7113386685615233   0.7617959604597195   0.9051870326095596   0.43226125301318014   0.08849255108511994   0.05433382624393325   0.8439689231393155   0.3283135580223374   0.1657473824759974   0.33070826520019225   0.883948658939038   0.8816588154510037   0.9892019896734191   0.7490467789005655   0.14566480406605997
0.4738530909445154   0.7924678011215851   0.504299948950372   0.28200667192514944   0.7935046214851728   0.5478842702094413   0.16801482601528628   0.12950230954828026   0.6323378166407805   0.8365456016479181   0.4062188655555667   0.2243152769387207   0.20007656362760032   0.7480530505627981   0.35188503931163345   0.3803463537994052   0.871763005605263   0.5823056680868007   0.021176774111441206   0.4963976948603672   0.9901041901542592   0.5931036784133817   0.2721299952108757   0.35073289079430725   0.5162510992097439   0.8006358772917966   0.7678300462605038   0.06872621886915782   0.7227464777245711   0.2527516070823552   0.5998152202452175   0.9392239093208775   0.09040866108379066   0.41620600543443714   0.19359635468965078   0.7149086323821569   0.8903320974561904   0.668152954871639   0.8417113153780174   0.3345622785827517   0.018569091850927394   0.08584728678483818   0.8205345412665761   0.8381645837223844   0.02846490169666813   0.4927436083714565   0.5484045460557003   0.48743169292807725   0.5122138024869243   0.6921077310796598   0.7805744997951966   0.41870547405891945   0.7894673247623532   0.4393561239973046   0.1807592795499791   0.4794815647380419   0.6990586636785625   0.023150118562867507   0.9871629248603283   0.764572932355885   0.8087265662223722   0.3549971636912286   0.14545160948231103   0.4300106537731333
0.7901574743714448   0.26914987690639036   0.3249170682157349   0.5918460700507487   0.7616925726747766   0.7764062685349339   0.7765125221600345   0.10441437712267153   0.2494787701878524   0.08429853745527403   0.995938022364838   0.6857089030637521   0.46001144542549927   0.6449424134579694   0.8151787428148588   0.20622733832571022   0.7609527817469368   0.6217922948951019   0.8280158179545305   0.4416544059698252   0.9522262155245647   0.2667951312038733   0.6825642084722194   0.011643752196691929   0.1620687411531199   0.997645254297483   0.3576471402564846   0.41979768214594315   0.4003761684783433   0.22123898576254902   0.58113461809645   0.3153833050232716   0.1508973982904909   0.136940448307275   0.5851965957316121   0.6296744019595195   0.6908859528649917   0.4919980348493056   0.7700178529167532   0.4234470636338093   0.9299331711180548   0.8702057399542037   0.9420020349622227   0.981792657663984   0.9777069555934902   0.6034106087503304   0.2594378264900032   0.9701489054672922   0.8156382144403703   0.6057653544528474   0.9017906862335187   0.550351223321349   0.41526204596202704   0.3845263686902984   0.32065606813706865   0.2349679182980774   0.26436464767153617   0.24758592038302338   0.7354594724054566   0.6052935163385579   0.5734786948065446   0.7555878855337178   0.9654416194887034   0.1818464527047486
0.6435455236884897   0.8853821455795141   0.023439584526480706   0.20005379504076454   0.6658385680949994   0.28197153682918374   0.7640017580364775   0.2299048895734724   0.8502003536546291   0.6762061823763363   0.8622110718029589   0.6795536662521234   0.43493830769260206   0.29167981368603796   0.5415550036658903   0.44458574795404604   0.17057366002106591   0.04409389330301459   0.8060955312604337   0.8392922316154882   0.5970949652145214   0.2885060077692968   0.8406539117717302   0.6574457789107395   0.9535494415260317   0.40312386218978274   0.8172143272452496   0.457391983869975   0.28771087343103224   0.121152325360599   0.05321256920877204   0.22748709429650255   0.4375105197764031   0.44494614298426266   0.19100149740581318   0.5479334280443792   0.002572212083801019   0.15326632929822473   0.6494464937399229   0.1033476800903331   0.8319985520627351   0.10917243599521013   0.8433509624794893   0.26405544847484497   0.23490358684821372   0.8206664282259133   0.002697050707759057   0.6066096695641054   0.281354145322182   0.4175425660361306   0.18548272346250952   0.1492176856941305   0.9936432718911498   0.2963902406755316   0.13227015425373748   0.9217305913976279   0.5561327521147467   0.8514440976912689   0.9412686568479243   0.3737971633532488   0.5535605400309457   0.6981777683930442   0.29182216310800135   0.27044948326291574
0.7215619879682106   0.589005332397834   0.44847120062851203   0.0063940347880707404   0.4866584011199968   0.7683389041719207   0.445774149920753   0.39978436522396527   0.2053042557978148   0.35079633813579014   0.2602914264582435   0.25056667952983475   0.21166098390666505   0.05440609746025855   0.128021272204506   0.3288360881322068   0.6555282317919183   0.2029619997689896   0.18675261535658172   0.955038924778958   0.1019676917609727   0.5047842313759454   0.8949304522485804   0.6845894415160423   0.3804057037927621   0.9157788989781113   0.44645925162006833   0.6781954067279715   0.8937473026727653   0.14743999480619055   0.0006851016993153572   0.27841104150400625   0.6884430468749505   0.7966436566704004   0.7403936752410719   0.027844361974171485   0.47678206296828546   0.7422375592101419   0.6123724030365659   0.6990082738419646   0.8212538311763671   0.5392755594411522   0.4256197876799842   0.7439693490630067   0.7192861394153944   0.034491328065206855   0.5306893354314038   0.0593799075469644   0.33888043562263226   0.11871242908709555   0.0842300838113355   0.38118450081899286   0.44513313294986695   0.971272434280905   0.08354498211202013   0.1027734593149866   0.7566900860749165   0.17462877761050458   0.34315130687094825   0.07492909734081513   0.279908023106631   0.4323912184003627   0.7307789038343824   0.3759208234988505
0.4586541919302639   0.8931156589592105   0.30515911615439817   0.6319514744358438   0.7393680525148695   0.8586243308940036   0.7744697807229943   0.5725715668888793   0.4004876168922373   0.739911901806908   0.6902396969116589   0.1913870660698865   0.9553544839423703   0.7686394675260031   0.6066947147996387   0.0886136067548999   0.19866439786745385   0.5940106899154985   0.26354340792869047   0.013684509414084785   0.9187563747608228   0.16161947151513578   0.5327645040943081   0.6377636859152344   0.4601021828305589   0.2685038125559253   0.22760538793990995   0.005812211479390542   0.7207341303156894   0.4098794816619217   0.45313560721691565   0.43324064459051115   0.3202465134234521   0.6699675798550137   0.7628959103052568   0.24185357852062464   0.36489202948108185   0.9013281123290106   0.1562011955056181   0.15323997176572474   0.166227631613628   0.307317422413512   0.8926577875769276   0.13955546235163996   0.24747125685280516   0.14569795089837623   0.3598932834826195   0.5017917764364056   0.7873690740222462   0.877194138342451   0.13228789554270956   0.49597956495701506   0.06663494370655683   0.46731465668052924   0.679152288325794   0.06273892036650393   0.7463884302831046   0.7973470768255156   0.9162563780205372   0.8208853418458792   0.38149640080202285   0.8960189644965051   0.7600551825149191   0.6676453700801546
0.21526876918839485   0.5887015420829931   0.8673973949379914   0.5280899077285146   0.9677975123355897   0.44300359118461685   0.5075041114553719   0.02629813129210897   0.1804284383133435   0.565809452842166   0.37521621591266235   0.5303185663350939   0.11379349460678664   0.09849479616163671   0.6960639275868684   0.46757964596859   0.367405064323682   0.30114771933612106   0.7798075495663312   0.6466943041227107   0.9859086635216591   0.40512875483961597   0.01975236705141217   0.9790489340425561   0.7706398943332643   0.8164272127566229   0.15235497211342072   0.45095902631404156   0.8028423819976745   0.373423621572006   0.6448508606580489   0.4246608950219326   0.6224139436843311   0.80761416872984   0.26963464474538645   0.8943423286868387   0.5086204490775444   0.7091193725682033   0.573570717158518   0.42676268271824874   0.14121538475386247   0.4079716532320823   0.7937631675921868   0.780068378595538   0.15530672123220335   0.0028428983924663025   0.7740108005407746   0.8010194445529819   0.3846668268989391   0.18641568563584343   0.6216558284273539   0.35006041823894035   0.5818244449012645   0.8129920640638374   0.9768049677693051   0.9253995232170078   0.9594105012169335   0.005377895333997361   0.7071703230239187   0.031057194530169065   0.45079005213938905   0.296258522765794   0.1335996058654006   0.6042945118119204
0.3095746673855266   0.8882868695337117   0.33983643827321375   0.8242261332163823   0.1542679461533232   0.8854439711412454   0.5658256377324391   0.023206688663400442   0.7696011192543841   0.699028285505402   0.9441698093050852   0.6731462704244601   0.1877766743531196   0.8860362214415646   0.9673648415357801   0.7477467472074524   0.22836617313618612   0.8806583261075672   0.26019451851186143   0.7166895526772833   0.7775761209967971   0.5843998033417732   0.12659491264646083   0.11239504086536295   0.46800145361127055   0.6961129338080615   0.7867584743732471   0.2881689076489806   0.3137335074579473   0.8106689626668161   0.22093283664080793   0.2649622189855802   0.5441323882035632   0.11164067716141404   0.2767630273357227   0.5918159485611201   0.3563557138504436   0.22560445571984947   0.30939818579994266   0.8440692013536677   0.1279895407142575   0.3449461296122822   0.04920366728808123   0.1273796486763844   0.3504134197174604   0.760546326270509   0.9226087546416204   0.014984607811021462   0.8824119661061899   0.06443339246244754   0.13585028026837334   0.7268157001620409   0.5686784586482425   0.2537644297956315   0.9149174436275654   0.46185348117646063   0.024546070444679307   0.14212375263421745   0.6381544162918427   0.8700375326153406   0.6681903565942356   0.916519296914368   0.3287562304919   0.025968331261672868
0.5402008158799781   0.5715731673020857   0.27955256320381877   0.8985886825852885   0.1897873961625178   0.8110268410315767   0.3569438085621984   0.883604074774267   0.30737543005632795   0.7465934485691291   0.22109352829382503   0.15678837461222617   0.7386969714080854   0.49282901877349766   0.3061760846662596   0.6949348934357655   0.7141509009634062   0.3507052661392802   0.668021668374417   0.824897360820425   0.04596054436917046   0.4341859692249122   0.33926543788251695   0.7989290295587521   0.5057597284891923   0.8626128019228264   0.0597128746786982   0.9003403469734637   0.31597233232667443   0.05158596089124973   0.7027690661164998   0.01673627219919661   0.008596902270346476   0.30499251232212055   0.4816755378226748   0.8599478975869704   0.269899930862261   0.8121634935486228   0.17549945315641519   0.16501300415120493   0.5557490298988549   0.46145822740934267   0.5074777847819982   0.34011564333078   0.5097884855296844   0.027272258184430444   0.16821234689948125   0.5411866137720279   0.004028757040492156   0.164659456261604   0.10849947222078306   0.6408462667985644   0.6880564247138177   0.11307349537035427   0.40573040610428324   0.6241099945993677   0.6794595224434712   0.8080809830482337   0.9240548682816084   0.7641620970123972   0.4095595915812102   0.9959174894996109   0.7485554151251932   0.5991490928611923
0.8538105616823554   0.5344592620902682   0.24107763034319502   0.2590334495304123   0.34402207615267094   0.5071870039058377   0.07286528344371375   0.7178468357583844   0.3399933191121788   0.34252754764423377   0.9643658112229306   0.07700056895982005   0.6519368943983611   0.2294540522738795   0.5586354051186475   0.4528905743604523   0.9724773719548898   0.42137306922564577   0.6345805368370391   0.6887284773480551   0.5629177803736796   0.4254555797260349   0.8860251217118458   0.08957938448686271   0.7091072186913243   0.8909963176357667   0.6449474913686508   0.8305459349564503   0.3650851425386533   0.383809313729929   0.572082207924937   0.11269909919806602   0.025091823426474574   0.04128176608569521   0.6077163967020064   0.03569853023824597   0.37315492902811354   0.8118277138118157   0.04908099158335893   0.5828079558777937   0.40067755707322367   0.39045464458616996   0.4145004547463199   0.8940794785297386   0.837759776699544   0.964999064860135   0.528475333034474   0.8045000940428759   0.1286525580082198   0.0740027472243683   0.8835278416658232   0.9739541590864255   0.7635674154695664   0.6901934334944393   0.3114456337408862   0.8612550598883595   0.7384755920430919   0.6489116674087441   0.7037292370388798   0.8255565296501135   0.36532066301497834   0.8370839535969284   0.6546482454555209   0.24274857377231984
0.9646431059417547   0.4466293090107584   0.24014779070920098   0.3486690952425813   0.1268833292422106   0.48163024415062344   0.7116724576747269   0.5441690011997053   0.9982307712339908   0.40762749692625516   0.8281446160089037   0.5702148421132799   0.23466335576442435   0.7174340634318158   0.5166989822680175   0.7089597822249204   0.4961877637213325   0.06852239602307171   0.8129697452291377   0.8834032525748069   0.1308671007063541   0.23143844242614334   0.15832149977361681   0.640654678802487   0.16622399476459943   0.7848091334153848   0.9181737090644159   0.29198558355990584   0.03934066552238882   0.30317888926476144   0.20650125138968892   0.7478165823602004   0.041109894288398   0.8955513923385063   0.37835663538078523   0.17760174024692055   0.8064465385239736   0.1781173289066905   0.8616576531127678   0.4686419580220001   0.3102587748026412   0.10959493288361877   0.048687907883630095   0.5852387054471931   0.17939167409628706   0.8781564904574755   0.8903664081100133   0.9445840266447061   0.013167679331687623   0.09334735704209056   0.9721926990455975   0.6525984430848003   0.9738270138092988   0.7901684677773291   0.7656914476559086   0.9047818607245998   0.9327171195209008   0.8946170754388229   0.38733481227512334   0.7271801204776792   0.12627058099692717   0.7164997465321323   0.5256771591623556   0.2585381624556792
0.816011806194286   0.6069048136485136   0.47698925127872543   0.673299457008486   0.636620132097999   0.7287483231910381   0.5866228431687122   0.72871543036378   0.6234524527663113   0.6354009661489476   0.6144301441231147   0.07611698727897966   0.6496254389570125   0.8452324983716184   0.8487386964672061   0.17133512655437985   0.7169083194361117   0.9506154229327957   0.4614038841920828   0.4441550060767006   0.5906377384391845   0.2341156764006633   0.9357267250297272   0.18561684362102143   0.7746259322448985   0.6272108627521498   0.45873747375100177   0.5123173866125355   0.13800580014689962   0.8984625395611116   0.8721146305822897   0.7836019562487555   0.5145533473805883   0.263061573412164   0.25768448645917497   0.7074849689697759   0.8649279084235758   0.41782907504054556   0.40894578999196884   0.536149842415396   0.14801958898746406   0.46721365210774995   0.9475419057998861   0.09199483633869542   0.5573818505482795   0.23309797570708665   0.011815180770158775   0.9063779927176739   0.782755918303381   0.6058871129549369   0.5530777070191569   0.3940606061051386   0.6447501181564813   0.7074245733938254   0.6809630764368674   0.6104586498563831   0.13019677077589306   0.4443629999816613   0.4232785899776924   0.9029736808866072   0.2652688623523173   0.026533924941115714   0.014332799985723578   0.3668238384712112
0.11724927336485325   0.5593202728333657   0.06679089418583756   0.2748290021325158   0.5598674228165738   0.3262222971262791   0.05497571341567878   0.3684510094148418   0.7771115045131928   0.7203351841713421   0.5018980063965218   0.9743904033097033   0.13236138635671146   0.012910610777516849   0.8209349299596544   0.3639317534533202   0.0021646155808183977   0.5685476107958556   0.39765633998196204   0.46095807256671295   0.7368957532285011   0.5420136858547399   0.38332353999623847   0.09413423409550174   0.6196464798636478   0.982693413021374   0.3165326458104009   0.819305231962986   0.05977905704707411   0.656471115895095   0.26155693239472216   0.45085422254814417   0.2826675525338813   0.9361359317237528   0.7596589259982004   0.4764638192384409   0.15030616617716985   0.923225320946236   0.9387239960385458   0.11253206578512075   0.14814155059635145   0.3546777101503804   0.5410676560565838   0.6515739932184078   0.4112457973678504   0.8126640242956406   0.15774411606034536   0.5574397591229061   0.7915993175042025   0.8299706112742665   0.8412114702499445   0.7381345271599201   0.7318202604571283   0.1734994953791715   0.5796545378552223   0.28728030461177595   0.4491527079232471   0.23736356365541872   0.819995611857022   0.8108164853733351   0.2988465417460772   0.3141382427091828   0.8812716158184761   0.6982844195882143
0.15070499114972574   0.9594605325588024   0.3402039597618922   0.04671042636980651   0.7394591937818754   0.14679650826316182   0.1824598437015469   0.48927066724690044   0.9478598762776729   0.31682589698889535   0.3412483734516024   0.7511361400869804   0.2160396158205445   0.14332640160972382   0.7615938355963802   0.46385583547520437   0.7668869078972974   0.9059628379543051   0.9415982237393582   0.6530393501018693   0.46804036615122024   0.5918245952451223   0.06032660792088209   0.954754930513655   0.31733537500149445   0.63236406268632   0.7201226481589899   0.9080445041438485   0.577876181219619   0.48556755442315813   0.537662804457443   0.418773836896948   0.6300163049419462   0.1687416574342628   0.19641443100584055   0.6676376968099677   0.4139766891214017   0.025415255824538987   0.43482059540946044   0.20378186133476334   0.6470897812241042   0.11945241787023388   0.49322237167010224   0.550742511232894   0.17904941507288402   0.5276278226251115   0.4328957637492202   0.5959875807192391   0.8617140400713895   0.8952637599387916   0.7127731155902303   0.6879430765753906   0.2838378588517705   0.4096962055156334   0.17511031113278733   0.26916923967844253   0.6538215539098243   0.24095454808137057   0.9786958801269467   0.6015315428684749   0.2398448647884226   0.21553929225683158   0.5438752847174864   0.39774968153371154
0.5927550835643184   0.09608687438659771   0.050652913047384104   0.8470071703008175   0.41370566849143436   0.5684590517614861   0.6177571492981639   0.2510195895815785   0.5519916284200448   0.6731952918226947   0.9049840337079337   0.5630765130061879   0.26815376956827436   0.26349908630706126   0.7298737225751463   0.29390727332774536   0.6143322156584501   0.022544538225690684   0.7511778424481995   0.6923757304592705   0.37448735087002744   0.8070052459688591   0.20730255773071316   0.294626048925559   0.7817322673057091   0.7109183715822613   0.15664964468332906   0.4476188786247415   0.36802659881427474   0.1424593198207752   0.5388924953851651   0.196599289043163   0.8160349703942299   0.4692640279980806   0.6339084616772315   0.6335227760369752   0.5478812008259556   0.2057649416910193   0.9040347391020852   0.33961550270922974   0.9335489851675055   0.1832204034653286   0.1528568966538857   0.6472397722499592   0.559061634297478   0.3762151574964695   0.9455543389231725   0.3526137233244002   0.777329366991769   0.6652967859142082   0.7889046942398434   0.9049948446996587   0.4093027681774942   0.522837466093433   0.25001219885467835   0.7083955556564957   0.5932677977832643   0.05357343809535236   0.6161037371774468   0.0748727796195206   0.045386596957308754   0.8478084964043331   0.7120689980753616   0.7352572769102909
0.11183761178980324   0.6645880929390044   0.559212101421476   0.08801750466033166   0.5527759774923252   0.2883729354425349   0.6136577624983035   0.7354037813359314   0.7754466105005562   0.6230761495283268   0.82475306825846   0.8304089366362727   0.36614384232306196   0.10023868343489385   0.5747408694037817   0.12201338097977701   0.7728760445397976   0.046665245339541486   0.9586371322263347   0.047140601360256426   0.7274894475824889   0.19885674893520844   0.24656813415097312   0.3118833244499656   0.6156518357926857   0.534268655996204   0.6873560327294971   0.2238658197896339   0.06287585830036045   0.24589572055366912   0.07369827023119366   0.48846203845370245   0.2874292477998043   0.6228195710253424   0.24894520197273365   0.6580531018174297   0.9212854054767423   0.5225808875904485   0.674204332568952   0.5360397208376527   0.14840936093694468   0.475915642250907   0.7155672003426172   0.4888991194773963   0.42091991335445583   0.27705889331569855   0.4689990661916441   0.17701579502743073   0.8052680775617702   0.7427902373194946   0.781643033462147   0.9531499752377969   0.7423922192614097   0.49689451676582547   0.7079447632309533   0.46468793678409437   0.45496297146160547   0.8740749457404831   0.45899956125821967   0.8066348349666647   0.5336775659848632   0.3514940581500346   0.7847952286892677   0.27059511412901194
0.3852682050479185   0.8755784158991277   0.06922802834665044   0.7816959946516157   0.9643482916934627   0.598519522583429   0.6002289621550063   0.6046801996241848   0.15908021413169246   0.8557292852639344   0.8185859286928594   0.6515302243863881   0.41668799487028274   0.358834768498109   0.11064116546190604   0.18684228760229368   0.9617250234086773   0.4847598227576259   0.6516416042036863   0.38020745263562905   0.42804745742381406   0.13326576460759132   0.8668463755144187   0.10961233850661713   0.04277925237589558   0.2576873487084637   0.7976183471677682   0.3279163438550015   0.07843096068243294   0.6591678261250347   0.19738938501276193   0.7232361442308166   0.9193507465507404   0.8034385408611002   0.3788034563199026   0.07170591984442856   0.5026627516804577   0.44460377236299115   0.26816229085799653   0.8848636322421349   0.5409377282717805   0.9598439496053652   0.6165206866543101   0.5046561796065059   0.11289027084796646   0.8265781849977739   0.7496743111398915   0.3950438410998887   0.07011101847207088   0.5688908362893101   0.9520559639721231   0.06712749724488719   0.991680057789638   0.9097230101642756   0.7546665789593612   0.3438913530140706   0.07232931123889748   0.10628446930317537   0.37586312263945865   0.272185433169642   0.5696665595584397   0.6616806969401843   0.1077008317814621   0.3873218009275071
0.028728831286659186   0.701836747334819   0.49118014512715197   0.8826656213210012   0.9158385604386927   0.8752585623370451   0.7415058339872606   0.4876217802211126   0.8457275419666218   0.30636772604773493   0.7894498700151373   0.4204942829762254   0.8540474841769838   0.3966447158834594   0.03478329105577614   0.07660292996215481   0.7817181729380864   0.29036024658028403   0.6589201684163175   0.8044174967925128   0.2120516133796467   0.6286795496400998   0.5512193366348555   0.41709569586500567   0.18332278209298752   0.9268428023052808   0.060039191507703454   0.5344300745440044   0.2674842216542948   0.051584239968235655   0.31853335752044293   0.046808294322891825   0.42175667968767294   0.7452165139205007   0.5290834875053055   0.6263140113466664   0.5677091955106891   0.34857179803704136   0.49430019644952944   0.5497110813845116   0.7859910225726027   0.058211551456757334   0.835380028033212   0.7452935845919988   0.5739394091929559   0.4295320018166575   0.28416069139835654   0.3281978887269931   0.3906166270999684   0.5026891995113768   0.22412149989065308   0.7937678141829887   0.12313240544567365   0.4511049595431411   0.9055881423702101   0.7469595198600969   0.7013757257580007   0.7058884456226404   0.37650465486490453   0.12064550851343046   0.13366653024731162   0.357316647585599   0.8822044584153751   0.5709344271289188
0.34767550767470895   0.2991050961288417   0.04682443038216315   0.82564084253692   0.7737360984817531   0.8695730943121841   0.7626637389838066   0.49744295380992687   0.3831194713817846   0.3668838948008074   0.5385422390931535   0.7036751396269382   0.25998706593611093   0.9157789352576663   0.6329540967229433   0.9567156197668412   0.5586113401781102   0.2098904896350259   0.2564494418580388   0.8360701112534108   0.42494480993079864   0.8525738420494269   0.3742449834426637   0.26513568412449195   0.07726930225608965   0.5534687459205851   0.32742055306050055   0.4394948415875719   0.3035332037743366   0.683895651608401   0.564756814076694   0.942051887777645   0.9204137323925521   0.31701175680759364   0.026214574983540444   0.23837674815070695   0.6604266664564411   0.40123282154992734   0.39326047826059707   0.28166112838386576   0.1018153262783309   0.19134233191490146   0.13681103640255826   0.44559101713045496   0.6768705163475323   0.3387684898654746   0.7625660529598945   0.18045533300596303   0.5996012140914426   0.7852997439448894   0.435145499899394   0.7409604914183912   0.296068010317106   0.10140409233648841   0.8703886858227   0.798908603640746   0.37565427792455397   0.7843923355288948   0.8441741108391596   0.560531855490039   0.7152276114681129   0.3831595139789674   0.4509136325785625   0.27887072710617333
0.6134122851897819   0.19181718206406595   0.3141025961760042   0.8332797099757184   0.9365417688422496   0.8530486921985914   0.5515365432161097   0.6528243769697554   0.336940554750807   0.06774894825370192   0.1163910433167157   0.9118638855513642   0.040872544433700954   0.9663448559172135   0.24600235749401567   0.1129552819106182   0.665218266509147   0.18195252038831874   0.40182824665485606   0.5524234264205791   0.9499906550410342   0.7987930064093514   0.9509146140762935   0.27355269931440573   0.3365783698512523   0.6069758243452854   0.6368120179002893   0.44027298933868736   0.4000366010090027   0.753927132146694   0.08527547468417963   0.787448612368932   0.06309604625819569   0.6861781838929921   0.9688844313674639   0.8755847268175678   0.022223501824494736   0.7198333279757786   0.7228820738734483   0.7626294449069496   0.3570052353153477   0.5378808075874598   0.3210538272185922   0.2102060184863705   0.40701458027431353   0.7390878011781086   0.37013921314229864   0.9366533191719647   0.07043621042306128   0.1321119768328231   0.7333271952420093   0.49638032983327735   0.6703996094140586   0.37818484468612906   0.6480517205578297   0.7089317174643454   0.6073035631558629   0.6920066607931369   0.6791672891903657   0.8333469906467775   0.5850800613313681   0.9721733328173583   0.9562852153169175   0.07071754573982791
0.22807482601602044   0.4342925252298985   0.6352313880983252   0.8605115272534575   0.8210602457417069   0.6952047240517899   0.26509217495602666   0.9238582080814927   0.7506240353186456   0.5630927472189668   0.5317649797140174   0.42747787824821537   0.08022442590458702   0.18490790253283776   0.8837132591561877   0.71854616078387   0.4729208627487241   0.4929012417397008   0.20454596996582192   0.8851991701370925   0.8878408014173559   0.5207279089223424   0.24826075464890443   0.8144816243972646   0.6597659754013354   0.08643538369244402   0.6130293665505792   0.9539700971438072   0.8387057296596285   0.39123065964065407   0.3479371915945525   0.030111889062314472   0.08808169434098292   0.8281379124216872   0.8161722118805352   0.6026340108140992   0.00785726843639591   0.6432300098888495   0.9324589527243475   0.884087850030229   0.5349364056876719   0.1503287681491487   0.7279129827585257   0.9988886798931366   0.6470956042703159   0.6296008592268062   0.47965222810962116   0.184407055495872   0.9873296288689805   0.5431654755343622   0.866622861559042   0.23043695835206482   0.14862389920935193   0.1519348158937081   0.5186856699644895   0.20032506928975033   0.060542204868369   0.32379690347202084   0.7025134580839543   0.5976910584756512   0.052684936431973084   0.6805668935831714   0.7700545053596067   0.7136032084454221
0.5177485307443013   0.5302381254340226   0.042141522601081165   0.7147145285522856   0.8706529264739853   0.9006372662072164   0.56248929449146   0.5303074730564136   0.8833232976050048   0.35747179067285423   0.695866432932418   0.2998705147043487   0.7346993983956529   0.20553697477914612   0.17718076296792848   0.0995454454145984   0.674157193527284   0.8817400713071253   0.47466730488397413   0.5018543869389471   0.6214722570953108   0.20117317772395396   0.7046127995243674   0.7882511784935251   0.10372372635100961   0.6709350522899313   0.6624712769232862   0.07353664994123953   0.23307079987702428   0.7702977860827149   0.09998198243182622   0.543229176884826   0.3497475022720194   0.4128259954098607   0.40411554949940826   0.24335866218047725   0.6150481038763664   0.20728902063071455   0.2269347865314798   0.14381321676587885   0.9408909103490825   0.32554894932358924   0.7522674816475057   0.6419588298269316   0.3194186532537716   0.12437577159963531   0.047654682123138274   0.8537076513334066   0.21569492690276199   0.453440719309704   0.38518340519985206   0.7801710013921671   0.9826241270257378   0.683142933226989   0.28520142276802585   0.23694182450734108   0.6328766247537183   0.27031693781712834   0.8810858732686175   0.9935831623268638   0.017828520877351876   0.06302791718641382   0.6541510867371377   0.849769945560985
0.0769376105282694   0.7374789678628245   0.9018836050896322   0.2078111157340533   0.7575189572744978   0.6131031962631892   0.8542289229664939   0.3541034644006467   0.5418240303717359   0.15966247695348526   0.4690455177666418   0.5739324630084797   0.5591999033459981   0.4765195437264962   0.18384409499861595   0.3369906385011386   0.9263232785922798   0.20620260590936784   0.3027582217299984   0.34340747617427475   0.9084947577149279   0.14317468872295402   0.6486071349928606   0.49363753061328974   0.8315571471866585   0.40569572086012945   0.7467235299032284   0.28582641487923643   0.07403818991216071   0.7925925245969402   0.8924946069367347   0.9317229504785897   0.5322141595404248   0.632930047643455   0.42344908917009283   0.35779048747011005   0.9730142561944267   0.15641050391695877   0.23960499417147688   0.020799848968971506   0.04669097760214695   0.950207898007591   0.9368467724414785   0.6773923727946968   0.13819621988721903   0.807033209284637   0.28823963744861786   0.18375484218140706   0.3066390727005605   0.40133748842450745   0.5415161075453894   0.8979284273021706   0.23260088278839977   0.6087449638275673   0.6490215006086548   0.9662054768235809   0.7003867232479749   0.9758149161841122   0.22557241143856194   0.6084149893534708   0.7273724670535481   0.8194044122671534   0.985967417267085   0.5876151403844994
0.6806814894514012   0.8691965142595625   0.049120644825606595   0.9102227675898026   0.5424852695641822   0.06216330497492558   0.7608810073769887   0.7264679254083956   0.23584619686362165   0.6608258165504182   0.21936489983159935   0.8285394981062248   0.003245314075221892   0.05208085272285091   0.5703433992229445   0.862334021282644   0.30285859082724703   0.07626593653873867   0.34477098778438264   0.25391903192917314   0.5754861237736989   0.2568615242715852   0.35880357051729755   0.6663038915446738   0.8948046343222977   0.3876650100120227   0.309682925691691   0.7560811239548713   0.3523193647581156   0.32550170503709713   0.5488019183147023   0.029613198546475726   0.11647316789449391   0.664675888486679   0.3294370184831029   0.20107370044025083   0.11322785381927203   0.6125950357638281   0.7590936192601583   0.33873967915760683   0.810369262992025   0.5363290992250894   0.4143226314757757   0.08482064722843373   0.23488313921832613   0.2794675749535042   0.055519060958478125   0.41851675568375996   0.3400785048960284   0.8918025649414815   0.7458361352667872   0.6624356317288886   0.9877591401379128   0.5663008599043844   0.19703421695208492   0.6328224331824129   0.8712859722434189   0.9016249714177054   0.8675971984689821   0.43174873274216213   0.7580581184241468   0.2890299356538773   0.10850357920882372   0.09300905358455527
0.9476888554321219   0.7527008364287879   0.6941809477330481   0.008188406356121544   0.7128057162137957   0.4732332614752837   0.6386618867745699   0.5896716506723616   0.3727272113177673   0.5814306965338022   0.8928257515077828   0.927236018943473   0.38496807117985454   0.015129836629417824   0.6957915345556978   0.29441358576105997   0.5136820989364356   0.11350486521171244   0.8281943360867158   0.8626648530188978   0.7556239805122887   0.8244749295578351   0.7196907568778921   0.7696557994343426   0.8079351250801668   0.07177409312904724   0.025509809144844   0.761467393078221   0.09512940886637115   0.5985408316537636   0.3868479223702741   0.17179574240585938   0.7224021975486038   0.017110135119961338   0.49402217086249134   0.24455972346238647   0.3374341263687493   0.001980298490543514   0.7982306363067936   0.9501461377013265   0.8237520274323137   0.888475433278831   0.9700363002200778   0.0874812846824287   0.06812804692002492   0.06400050372099594   0.25034554334218573   0.3178254852480862   0.26019292183985804   0.9922264105919487   0.22483573419734174   0.5563580921698652   0.16506351297348687   0.3936855789381852   0.8379878118270676   0.3845623497640058   0.4426613154248831   0.37657544381822383   0.34396564096457627   0.1400026263016193   0.10522718905613376   0.3745951453276803   0.5457350046577828   0.18985648860029278
0.2814751616238201   0.48611971204884924   0.575698704437705   0.10237520391786407   0.2133471147037952   0.42211920832785327   0.32535316109551926   0.784549718669778   0.9531541928639372   0.4298927977359046   0.10051742689817754   0.22819162649991276   0.7880906798904503   0.036207218797719425   0.2625296150711099   0.8436292767359069   0.34542936446556727   0.6596317749794957   0.9185639741065336   0.7036266504342876   0.2402021754094335   0.2850366296518153   0.3728289694487508   0.5137701618339949   0.9587270137856134   0.798916917602966   0.7971302650110459   0.4113949579161308   0.7453798990818182   0.37679770927511275   0.4717771039155266   0.6268452392463529   0.792225706217881   0.9469049115392082   0.3712596770173491   0.3986536127464402   0.004135026327430726   0.9106976927414887   0.10873006194623916   0.5550243360105331   0.6587056618618634   0.25106591776199316   0.19016608783970554   0.8513976855762455   0.41850348645242996   0.9660292881101779   0.8173371183909547   0.33762752374225063   0.4597764726668166   0.1671123705072118   0.02020685337990884   0.9262325658261198   0.7143965735849984   0.790314661232099   0.5484297494643823   0.2993873265797669   0.9221708673671173   0.8434097496928908   0.1771700724470332   0.9007337138333268   0.9180358410396866   0.9327120569514021   0.06844001050079404   0.3457093778227936
0.25933017917782314   0.681646139189409   0.8782739226610885   0.4943116922465481   0.8408266927253931   0.7156168510792311   0.060936804270133794   0.15668416850429745   0.3810502200585766   0.5485044805720193   0.04072995089022496   0.23045160267817766   0.6666536464735783   0.7581898193399202   0.4923002014258427   0.9310642760984107   0.7444827791064609   0.9147800696470294   0.31513012897880954   0.030330562265084   0.8264469380667743   0.9820680126956273   0.24669011847801547   0.6846211844422905   0.5671167588889512   0.30042187350621835   0.368416195816927   0.19030949219574236   0.726290066163558   0.5848050224269873   0.3074793915467932   0.033625323691444914   0.3452398461049814   0.03630054185496801   0.26674944065656825   0.8031737210132672   0.6785861996314032   0.27811072251504776   0.7744492392307255   0.8721094449148565   0.9341034205249422   0.36333065286801836   0.459319110251916   0.8417788826497725   0.10765648245816796   0.38126264017239103   0.21262899177390054   0.1571576982074821   0.5405397235692168   0.08084076666617265   0.8442127959569735   0.9668482060117397   0.8142496574056588   0.49603574423918534   0.5367334044101804   0.9332228823202948   0.4690098113006774   0.45973520238421733   0.2699839637536121   0.13004916130702757   0.7904236116692742   0.1816244798691696   0.4955347245228866   0.25793971639217106
0.856320191144332   0.8182938270011513   0.03621561427097058   0.4161608337423985   0.748663708686164   0.4370311868287602   0.82358662249707   0.25900313553491644   0.20812398511694724   0.35619042016258756   0.9793738265400965   0.2921549295231767   0.39387432771128844   0.8601546759234022   0.4426404221299161   0.35893204720288185   0.924864516410611   0.40041947353918483   0.172656458376304   0.22888288589585432   0.13444090474133674   0.21879499367001526   0.6771217338534175   0.9709431695036833   0.27812071359700474   0.40050116666886404   0.6409061195824468   0.5547823357612848   0.5294570049108407   0.9634699798401039   0.8173194970853768   0.29577920022636833   0.3213330197938935   0.6072795596775162   0.8379456705452804   0.003624270703191666   0.9274586920826051   0.747124883754114   0.3953052484153642   0.6446922235003099   0.0025941756719940565   0.3467054102149292   0.22264879003906016   0.4158093376044555   0.8681532709306573   0.12791041654491392   0.5455270561856428   0.44486616810077223   0.5900325573336526   0.7274092498760499   0.9046209366031959   0.8900838323394875   0.06057555242281182   0.7639392700359461   0.0873014395178191   0.5943046321131191   0.7392425326289184   0.15665971035842985   0.2493557689725388   0.5906803614099274   0.8117838405463133   0.4095348266043158   0.8540505205571747   0.9459881379096177
0.8091896648743192   0.06282941638938662   0.6314017305181144   0.5301788003051622   0.9410363939436619   0.9349189998444727   0.08587467433247173   0.08531263220438992   0.35100383661000933   0.20750974996842278   0.18125373772927583   0.19522879986490246   0.2904282841871975   0.44357047993247667   0.09395229821145673   0.6009241677517834   0.5511857515582792   0.2869107695740468   0.8445965292389179   0.010243806341855897   0.739401911011966   0.877375942969731   0.9905460086817433   0.06425566843223826   0.9302122461376467   0.8145465265803444   0.3591442781636288   0.5340768681270761   0.9891758521939849   0.8796275267358717   0.2732696038311571   0.4487642359226862   0.6381720155839755   0.6721177767674489   0.09201586610188126   0.2535354360577837   0.34774373139677794   0.22854729683497227   0.9980635678904245   0.6526112683060004   0.7965579798384987   0.9416365272609254   0.1534670386515066   0.6423674619641445   0.05715606882653277   0.06426058429119444   0.1629210299697633   0.5781117935319062   0.12694382268888604   0.24971405771085003   0.8037767518061345   0.04403492540483012   0.1377679704949012   0.37008653097497834   0.5305071479749773   0.5952706894821439   0.49959595491092573   0.6979687542075294   0.4384912818730961   0.3417352534243602   0.1518522235141478   0.46942145737255714   0.4404277139826716   0.6891239851183598
0.3552942436756491   0.5277849301116317   0.286960675331165   0.04675652315421532   0.2981381748491163   0.4635243458204373   0.12403964536140172   0.4686447296223091   0.17119435216023027   0.21381028810958722   0.32026289355526727   0.42460980421747896   0.03342638166532908   0.8437237571346089   0.7897557455802899   0.8293391147353351   0.5338304267544034   0.1457550029270795   0.3512644637071938   0.48760386131097483   0.38197820324025555   0.6763335455545223   0.9108367497245222   0.7984798761926151   0.02668395956460647   0.14854861544289066   0.6238760743933572   0.7517233530383997   0.7285457847154901   0.6850242696224534   0.49983642903195546   0.2830786234160906   0.5573514325552599   0.4712139815128662   0.17957353547668822   0.8584688191986116   0.5239250508899308   0.6274902243782573   0.3898177898963983   0.0291297044632766   0.9900946241355274   0.4817352214511778   0.038553326189204554   0.5415258431523018   0.6081164208952718   0.8054016758966555   0.12771657646468237   0.7430459669596867   0.5814324613306654   0.6568530604537648   0.5038405020713251   0.9913226139212871   0.8528866766151753   0.9718287908313115   0.0040040730393697   0.7082439905051965   0.2955352440599154   0.5006148093184453   0.8244305375626815   0.8497751713065848   0.7716101931699846   0.873124584940188   0.43461274766628316   0.8206454668433082
0.7815155690344572   0.39138936348901016   0.39605942147707857   0.27911962369100646   0.17339914813918525   0.5859876875923546   0.2683428450123962   0.5360736567313197   0.5919666868085198   0.9291346271385899   0.764502342941071   0.5447510428100326   0.7390800101933446   0.9573058363072785   0.7604982699017013   0.8365070523048362   0.4435447661334292   0.45669102698883324   0.9360677323390199   0.9867318809982514   0.6719345729634446   0.5835664420486453   0.5014549846727367   0.16608641415494318   0.8904190039289874   0.19217707855963517   0.10539556319565814   0.8869667904639368   0.7170198557898022   0.6061893909672805   0.8370527181832619   0.35089313373261705   0.12505316898128235   0.6770547638286907   0.07255037524219088   0.8061420909225844   0.3859731587879378   0.7197489275214122   0.31205210534048955   0.9696350386177481   0.9424283926545086   0.26305790053257894   0.37598437300146964   0.9829031576194968   0.270493819691064   0.6794914584839337   0.874529388328733   0.8168167434645536   0.3800748157620766   0.4873143799242985   0.7691338251330748   0.9298499530006168   0.6630549599722744   0.881124988957018   0.9320811069498129   0.5789568192679998   0.5380017909909921   0.20407022512832737   0.8595307317076221   0.7728147283454154   0.15202863220305426   0.48432129760691517   0.5474786263671325   0.8031796897276672
0.20960023954854567   0.22126339707433626   0.17149425336566282   0.8202765321081704   0.9391064198574817   0.5417719385904026   0.29696486503692987   0.003459788643616857   0.5590316040954051   0.05445755866610414   0.527831039903855   0.07360983564300001   0.8959766441231306   0.17333256970908614   0.5957499329540422   0.4946530163750002   0.3579748531321386   0.9692623445807588   0.7362192012464202   0.7218382880295848   0.20594622092908432   0.4849410469738436   0.18874057487928766   0.9186585983019175   0.9963459813805386   0.2636776498995073   0.01724632151362485   0.09838206619374713   0.05723956152305701   0.7219057113091047   0.720281456476695   0.09492227755013027   0.49820795742765195   0.6674481526430006   0.19245041657283993   0.021312441907130258   0.6022313133045213   0.49411558293391444   0.5967004836187978   0.5266594255321301   0.2442564601723827   0.5248532383531557   0.8604812823723776   0.8048211375025452   0.0383102392432984   0.03991219137931205   0.6717407074930899   0.8861625392006277   0.04196425786275974   0.7762345414798048   0.6544943859794651   0.7877804730068806   0.9847246963397027   0.05432883017069998   0.9342129295027701   0.6928581954567503   0.4865167389120508   0.3868806775276994   0.7417625129299302   0.67154575354962   0.8842854256075294   0.892765094593785   0.14506202931113243   0.14488632801748996
0.6400289654351468   0.3679118562406293   0.28458074693875485   0.3400651905149447   0.6017187261918484   0.32799966486131726   0.6128400394456649   0.45390265131431706   0.5597544683290886   0.5517651233815125   0.9583456534661998   0.6661221783074365   0.5750297719893859   0.49743629321081256   0.02413272396342975   0.9732639828506863   0.0885130330773351   0.1105556156831132   0.2823702110334996   0.30171822930106623   0.20422760746980562   0.21779052108932825   0.13730818172236714   0.15683190128357627   0.5641986420346589   0.8498786648486989   0.8527274347836123   0.8167667107686315   0.9624799158428105   0.5218789999873817   0.23988739533794737   0.3628640594543145   0.40272544751372186   0.9701138766058691   0.2815417418717475   0.696741881146878   0.827695675524336   0.47267758339505656   0.25740901790831777   0.7234778982961917   0.7391826424470008   0.3621219677119434   0.9750388068748183   0.42175966899512546   0.5349550349771952   0.14433144662261513   0.8377306251524511   0.2649277677115492   0.9707563929425364   0.29445278177391615   0.9850031903688388   0.44816105694291763   0.00827647709972592   0.7725737817865345   0.7451157950308914   0.08529699748860317   0.605551029586004   0.8024599051806653   0.46357405315914385   0.3885551163417252   0.7778553540616681   0.3297823217856088   0.20616503525082608   0.6650772180455334
0.03867271161466722   0.9676603540736654   0.23112622837600788   0.243317549050408   0.5037176766374719   0.8233289074510503   0.3933956032235568   0.9783897813388588   0.5329612836949356   0.528876125677134   0.40839241285471806   0.5302287243959412   0.5246848065952097   0.7563023438905996   0.6632766178238266   0.44493172690733795   0.9191337770092056   0.9538424387099343   0.19970256466468278   0.056376610565612766   0.1412784229475375   0.6240601169243255   0.9935375294138566   0.3912993925200793   0.10260571133287028   0.6563997628506602   0.7624113010378488   0.14798184346967128   0.5988880346953983   0.8330708553996099   0.369015697814292   0.16959206213081246   0.06592675100046275   0.30419472972247574   0.9606232849595739   0.6393633377348713   0.5412419444052531   0.5478923858318762   0.2973466671357473   0.19443161082753335   0.6221081673960475   0.5940499471219418   0.09764410247106453   0.1380550002619206   0.48082974444851   0.9699898301976163   0.10410657305720784   0.7467556077418414   0.37822403311563974   0.31359006734695616   0.341695272019359   0.59877376427217   0.7793359984202415   0.4805192119473463   0.972679574205067   0.4291817021413576   0.7134092474197787   0.17632448222487054   0.012056289245493072   0.7898183644064862   0.17216730301452557   0.6284320963929945   0.7147096221097458   0.5953867535789529
0.5500591356184781   0.03438214927105256   0.6170655196386813   0.4573317533170323   0.06922939116996804   0.06439231907343625   0.5129589465814733   0.710576145575191   0.6910053580543283   0.7508022517264801   0.17126367456211436   0.11180238130302092   0.9116693596340869   0.27028303977913376   0.19858410035704735   0.6826206791616634   0.1982601122143082   0.09395855755426319   0.18652781111155425   0.8928023147551771   0.02609280919978261   0.4655264611612688   0.4718181890018085   0.2974155611762242   0.47603367358130455   0.43114431189021624   0.8547526693631273   0.8400838078591919   0.4068042824113365   0.36675199281677995   0.3417937227816539   0.12950766228400093   0.7157989243570082   0.6159497410902999   0.17053004821953952   0.017705280980980013   0.8041295647229213   0.34566670131116617   0.9719459478624922   0.33508460181931665   0.6058694525086131   0.251708143756903   0.785418136750938   0.4422822870641396   0.5797766433088305   0.7861816825956341   0.3135999477491294   0.14486672588791538   0.10374296972752597   0.35503737070541797   0.45884727838600214   0.3047829180287235   0.6969386873161895   0.988285377888638   0.11705355560434824   0.17527525574472255   0.9811397629591813   0.3723356367983381   0.9465235073848087   0.15756997476374254   0.17701019823625996   0.026668935487171922   0.9745775595223165   0.8224853729444258
0.5711407457276468   0.774960791730269   0.18915942277137862   0.3802030858802863   0.9913641024188163   0.9887791091346347   0.8755594750222492   0.2353363599923709   0.8876211326912904   0.6337417384292168   0.4167121966362471   0.9305534419636474   0.19068244537510087   0.6454563605405788   0.2996586410318988   0.7552781862189248   0.20954268241591958   0.2731207237422407   0.3531351336470901   0.5977082114551824   0.032532484179659614   0.2464517882550688   0.3785575741247736   0.7752228385107565   0.46139173845201276   0.47149099652479987   0.18939815135339494   0.3950197526304702   0.4700276360331964   0.4827118873901651   0.3138386763311457   0.1596833926380993   0.5824065033419061   0.8489701489609482   0.8971264796948986   0.22912995067445188   0.3917240579668052   0.20351378842036946   0.5974678386629998   0.473851764455527   0.18218137555088562   0.9303930646781288   0.24433270501590965   0.8761435530003447   0.14964889137122603   0.6839412764230599   0.8657751308911361   0.10092071448958821   0.6882571529192133   0.21245027989826012   0.6763769795377411   0.705900961859118   0.2182295168860168   0.729738392508095   0.36253830320659547   0.5462175692210187   0.6358230135441107   0.8807682435471468   0.46541182351169685   0.3170876185465668   0.24409895557730552   0.6772544551267773   0.8679439848486971   0.8432358540910397
0.06191758002641989   0.7468613904486485   0.6236112798327874   0.9670923010906951   0.9122686886551938   0.06292011402558857   0.7578361489416513   0.8661715866011068   0.22401153573598062   0.8504698341273285   0.08145916940391018   0.16027062474198886   0.005782018849963812   0.12073144161923341   0.7189208661973148   0.6140530555209701   0.3699590053058531   0.23996319807208666   0.25350904268561786   0.29696543697440336   0.12586004972854756   0.5627087429453094   0.3855650578369208   0.45372958288336357   0.06394246970212768   0.8158473524966608   0.7619537780041333   0.48663728179266846   0.1516737810469338   0.7529272384710722   0.00411762906248205   0.6204656951915616   0.9276622453109532   0.9024574043437438   0.9226584596585719   0.4601950704495727   0.9218802264609893   0.7817259627245104   0.20373759346125714   0.8461420149286025   0.5519212211551363   0.5417627646524238   0.9502285507756393   0.5491765779541993   0.4260611714265887   0.9790540217071144   0.5646634929387184   0.09544699507083566   0.36211870172446103   0.16320666921045357   0.8027097149345851   0.6088097132781672   0.21044492067752724   0.41027943073938133   0.7985920858721031   0.9883440180866057   0.28278267536657403   0.5078220263956374   0.8759336262135311   0.5281489476370329   0.3609024489055847   0.7260960636711271   0.672196032752274   0.6820069327084304
0.8089812277504485   0.18433329901870335   0.7219674819766347   0.13283035475423113   0.38292005632385967   0.20527927731158896   0.1573039890379163   0.037383359683395456   0.020801354599398643   0.0420726081011354   0.3545942741033312   0.42857364640522827   0.8103564339218714   0.6317931773617541   0.5560021882312282   0.4402296283186226   0.5275737585552973   0.12397115096611659   0.680068562017697   0.9120806806815898   0.1666713096497127   0.3978750872949895   0.00787252926542305   0.23007374797315938   0.35769008189926427   0.21354178827628612   0.2859050472887883   0.09724339321892825   0.9747700255754046   0.008262510964697154   0.12860105825087204   0.05986003353553279   0.9539686709760059   0.9661899028635618   0.7740067841475409   0.6312863871303045   0.14361223705413453   0.33439672550180766   0.21800459591631263   0.19105675881168194   0.6160384784988372   0.21042557453569105   0.5379360338986156   0.27897607813009223   0.44936716884912453   0.8125504872407016   0.5300635046331925   0.04890233015693284   0.09167708694986022   0.5990086989644154   0.24415845734440422   0.9516589369380046   0.11690706137445563   0.5907461879997183   0.11555739909353219   0.8917989034024718   0.16293839039844968   0.6245562851361566   0.34155061494599137   0.26051251627216726   0.019326153344315134   0.2901595596343489   0.12354601902967872   0.06945575746048532
0.40328767484547795   0.07973398509865784   0.5856099851310631   0.7904796793303931   0.9539205059963535   0.26718349785795625   0.055546480497870615   0.7415773491734603   0.8622434190464933   0.6681747988935408   0.8113880231534664   0.7899184122354557   0.7453363576720375   0.07742861089382254   0.6958306240599342   0.8981195088329839   0.582397967273588   0.452872325757666   0.35428000911394286   0.6376069925608167   0.5630718139292727   0.1627127661233171   0.23073399008426412   0.5681512351003313   0.15978413908379482   0.08297878102465926   0.645124004953201   0.7776715557699382   0.20586363308744138   0.815795283166703   0.5895775244553304   0.03609420659647791   0.34362021404094817   0.14762048427316216   0.7781895013018639   0.24617579436102224   0.5982838563689106   0.07019187337933963   0.08235887724192976   0.34805628552803836   0.015885889095322656   0.6173195476216736   0.728078868127987   0.7104492929672218   0.4528140751660499   0.45460678149835654   0.4973448780437228   0.14229805786689048   0.293029936082255   0.37162800047369726   0.8522208730905219   0.3646265020969523   0.08716630299481365   0.5558327173069942   0.26264334863519145   0.3285322955004744   0.7435460889538655   0.40821223303383214   0.4844538473333275   0.08235650113945214   0.1452622325849549   0.3380203596544925   0.4020949700913978   0.7343002156114138
0.12937634348963226   0.7207008120328189   0.6740161019634109   0.023850922644191988   0.6765622683235823   0.26609403053446234   0.17667122391968804   0.8815528647773015   0.3835323322413273   0.8944660300607651   0.32445035082916623   0.5169263626803492   0.2963660292465137   0.3386333127537708   0.06180700219397474   0.1883940671798748   0.5528199402926482   0.9304210797199387   0.5773531548606472   0.10603756604042268   0.4075577077076933   0.5924007200654462   0.17525818476924948   0.3717373504290089   0.27818136421806106   0.8716999080326273   0.5012420828058386   0.34788642778481693   0.6016190958944786   0.605605877498165   0.3245708588861506   0.46633356300751544   0.2180867636531513   0.7111398474374   0.00012050805698439384   0.9494072003271662   0.9217207344066376   0.37250653468362915   0.9383135058630097   0.7610131331472914   0.3689007941139894   0.4420854549636905   0.36096035100236246   0.6549755671068688   0.9613430864062961   0.8496847348982444   0.18570216623311295   0.2832382166778598   0.683161722188235   0.977984826865617   0.6844600834272743   0.9353517888930428   0.0815426262937564   0.37237894936745203   0.3598892245411237   0.46901822588552744   0.8634558626406051   0.6612391019300521   0.35976871648413933   0.5196110255583613   0.9417351282339675   0.2887325672464229   0.4214552106211297   0.7585978924110698
0.5728343341199781   0.8466471122827324   0.06049485961876723   0.1036223253042011   0.611491247713682   0.996962377384488   0.8747926933856542   0.8203841086263413   0.928329525525447   0.018977550518871025   0.19033260995837997   0.8850323197332984   0.8467868992316906   0.646598601151419   0.8304433854172563   0.416014093847771   0.9833310365910855   0.985359499221367   0.47067466893311694   0.8964030682894097   0.04159590835711795   0.6966269319749441   0.04921945831198728   0.13780517587833993   0.4687615742371398   0.8499798196922117   0.98872459869322   0.03418285057413885   0.8572703265234578   0.8530174423077237   0.11393190530756578   0.21379874194779755   0.9289408009980108   0.8340398917888526   0.9235992953491858   0.32876642221449914   0.08215390176632024   0.18744129063743362   0.09315590993192957   0.9127523283667281   0.09882286517523478   0.20208179141606666   0.6224812409988126   0.016349260077318396   0.057226956818116834   0.5054548594411226   0.5732617826868254   0.8785440841989784   0.588465382580977   0.6554750397489109   0.5845371839936053   0.8443612336248396   0.7311950560575192   0.8024575974411873   0.4706052786860395   0.630562491677042   0.8022542550595084   0.9684177056523346   0.5470059833368537   0.30179606946254295   0.7201003532931882   0.780976415014901   0.45385007340492417   0.3890437410958148
0.6212774881179534   0.5788946235988343   0.8313688324061115   0.3726944810184964   0.5640505312998365   0.07343976415771172   0.25810704971928616   0.4941503968195179   0.9755851487188595   0.41796472440880084   0.6735698657256809   0.6497891631946783   0.24439009266134032   0.6155071269676136   0.20296458703964132   0.019226671517636244   0.4421358376018319   0.647089421315279   0.6559586037027876   0.7174306020550933   0.7220354843086437   0.866113006300378   0.20210853029786344   0.32838686095927855   0.10075799619069034   0.2872183827015437   0.37073969789175193   0.9556923799407822   0.5367074648908537   0.21377861854383198   0.11263264817246575   0.46154198312126427   0.5611223161719943   0.7958138941350311   0.4390627824467849   0.811752819926586   0.31673222351065394   0.1803067671674176   0.23609819540714358   0.7925261484089497   0.874596385908822   0.5332173458521385   0.580139591704356   0.07509554635385639   0.15256090160017832   0.6671043395517605   0.37803106140649256   0.7467086853945778   0.05180290540948797   0.3798859568502168   0.007291363514740645   0.7910163054537956   0.5150954405186342   0.16610733830638483   0.8946587153422749   0.32947432233253143   0.95397312434664   0.3702934441713537   0.45559593289549   0.5177215024059455   0.6372409008359861   0.1899866770039361   0.2194977374883464   0.7251953539969958
0.762644514927164   0.6567693311517975   0.6393581457839904   0.6500998076431393   0.6100836133269857   0.989664991600037   0.26132708437749785   0.9033911222485616   0.5582807079174977   0.6097790347498201   0.25403572086275716   0.11237481679476585   0.043185267398863504   0.4436716964434353   0.3593770055204823   0.7829004944622344   0.08921214305222357   0.07337825227208163   0.9037810726249923   0.265178992056289   0.4519712422162376   0.8833915752681455   0.684283335136646   0.5399836380592932   0.6893267272890736   0.22662224411634802   0.04492518935265553   0.8898838304161538   0.07924311396208793   0.23695725251631106   0.7835981049751577   0.9864927081675923   0.5209624060445902   0.627178217766491   0.5295623841124005   0.8741178913728265   0.47777713864572674   0.18350652132305564   0.17018537859191823   0.09121739691059202   0.38856499559350316   0.110128269050974   0.26640430596692594   0.826038404854303   0.9365937533772656   0.22673669378282846   0.58212097083028   0.28605476679500985   0.24726702608819204   0.00011444966648043158   0.5371957814776245   0.39617093637885603   0.1680239121261041   0.7631571971501694   0.7535976765024668   0.4096782282112637   0.6470615060815138   0.13597897938367845   0.22403529239006625   0.5355603368384373   0.16928436743578712   0.9524724580606229   0.05384991379814804   0.44434293992784524
0.7807193718422839   0.8423441890096488   0.7874456078312221   0.6183045350735422   0.8441256184650183   0.6156074952268203   0.20532463700094214   0.3322497682785323   0.5968585923768263   0.6154930455603399   0.6681288555233177   0.9360788318996763   0.4288346802507222   0.8523358484101705   0.9145311790208509   0.5264006036884126   0.7817731741692083   0.7163568690264921   0.6904958866307846   0.9908402668499753   0.6124888067334212   0.7638844109658693   0.6366459728326366   0.54649732692213   0.8317694348911373   0.9215402219562205   0.8492003650014145   0.9281927918485878   0.987643816426119   0.30593272672940014   0.6438757280004723   0.5959430235700556   0.3907852240492927   0.6904396811690602   0.9757468724771546   0.6598641916703792   0.9619505437985705   0.8381038327588897   0.06121569345630379   0.1334635879819667   0.18017736962936215   0.12174696373239756   0.37071980682551914   0.1426233211319914   0.5676885628959409   0.35786255276652823   0.7340738339928826   0.5961259942098613   0.7359191280048036   0.43632233081030775   0.8848734689914681   0.6679332023612735   0.7482753115786847   0.13038960408090763   0.24099774099099577   0.07199017879121794   0.35749008752939193   0.4399499229118474   0.2652508685138411   0.4121259871208387   0.3955395437308214   0.6018460901529578   0.20403517505753732   0.278662399138872
0.21536217410145925   0.48009912642056024   0.8333153682320181   0.1360390780068806   0.6476736112055184   0.12223657365403195   0.09924153423913558   0.5399130837970193   0.9117544832007147   0.6859142428437242   0.21436806524766747   0.8719798814357458   0.16347917162203016   0.5555246387628165   0.9733703242566717   0.7999897026445278   0.8059890840926383   0.11557471585096912   0.7081194557428306   0.38786371552368915   0.4104495403618168   0.5137286256980114   0.5040842806852933   0.10920131638481717   0.19508736626035755   0.03362949927745114   0.6707689124532751   0.9731622383779366   0.5474137550548392   0.9113929256234192   0.5715273782141396   0.43324915458091734   0.6356592718541244   0.225478682779695   0.3571593129664721   0.5612692731451716   0.47218010023209434   0.6699540440168784   0.3837889887098004   0.7612795705006438   0.6661910161394561   0.5543793281659093   0.6756695329669699   0.37341585497695456   0.2557414757776393   0.040650702467897974   0.17158525228167654   0.2642145385921374   0.06065410951728169   0.007021203190446834   0.5008163398284015   0.29105230021420087   0.5132403544624424   0.09562827756702766   0.9292889616142619   0.8578031456332835   0.877581082608318   0.8701495947873327   0.5721296486477897   0.29653387248811197   0.4054009823762237   0.20019555077045423   0.18834065993798935   0.5352543019874683
0.7392099662367676   0.6458162226045449   0.5126711269710196   0.16183844701051364   0.4834684904591284   0.6051655201366469   0.341085874689343   0.8976239084183762   0.42281438094184665   0.5981443169462001   0.8402695348609416   0.6065716082041754   0.9095740264794042   0.5025160393791724   0.9109805732466797   0.7487684625708919   0.031992943871086185   0.6323664445918398   0.33885092459889   0.45223459008277994   0.6265919614948625   0.43217089382138557   0.15051026466090064   0.9169802880953117   0.8873819952580949   0.7863546712168407   0.6378391376898811   0.7551418410847981   0.40391350479896654   0.18118915108019373   0.2967532630005381   0.8575179326664218   0.9810991238571198   0.5830448341339937   0.45648372813959653   0.25094632446224646   0.07152509737771565   0.0805287947548212   0.5455031548929168   0.5021778618913546   0.03953215350662946   0.44816235016298145   0.20665223029402682   0.04994327180857466   0.41294019201176696   0.015991456341595878   0.0561419656331262   0.13296298371326296   0.5255581967536721   0.22963678512475522   0.4183028279432451   0.3778211426284649   0.12164469195470559   0.04844763404456149   0.12154956494270697   0.520303209962043   0.14054556809758575   0.4654027999105679   0.6650658368031104   0.2693568854997966   0.0690204707198701   0.38487400515574666   0.11956268191019362   0.767179023608442
0.02948831721324063   0.9367116549927652   0.9129104516161668   0.7172357517998673   0.6165481252014736   0.9207201986511694   0.8567684859830406   0.5842727680866043   0.09098992844780156   0.6910834135264141   0.4384656580397955   0.20645162545813947   0.969345236493096   0.6426357794818526   0.3169160930970885   0.6861484154960964   0.8287996683955102   0.17723297957128478   0.6518502562939781   0.41679152999629987   0.7597791976756402   0.7923589744155382   0.5322875743837845   0.6496125063878578   0.7302908804623995   0.855647319422773   0.6193771227676177   0.9323767545879905   0.11374275526092584   0.9349271207716036   0.7626086367845771   0.3481039865013862   0.02275282681312429   0.24384370724518947   0.3241429787447816   0.1416523610432467   0.05340759032002833   0.6012079277633369   0.007226885647693077   0.4555039455471503   0.22460792192451812   0.42397494819205206   0.355376629353715   0.038712415550850414   0.464828724248878   0.6316159737765139   0.8230890549699306   0.38909990916299253   0.7345378437864785   0.775968654353741   0.20371193220231282   0.456723154575002   0.6207950885255527   0.8410415335821374   0.44110329541773574   0.10861916807361584   0.5980422617124284   0.597197826336948   0.11696031667295413   0.9669668070303691   0.5446346713924001   0.9959898985736111   0.10973343102526105   0.5114628614832188
0.3200267494678819   0.572014950381559   0.7543568016715461   0.4727504459323685   0.8551980252190039   0.9403989766050451   0.9312677467016156   0.08365053676937591   0.12066018143252547   0.16443032225130413   0.7275558144993027   0.6269273821943739   0.49986509290697284   0.3233887886691667   0.286452519081567   0.5183082141207581   0.9018228311945444   0.7261909623322187   0.16949220240861287   0.5513414070903889   0.35718815980214447   0.7302010637586076   0.059758771383351804   0.039878545607170066   0.03716141033426253   0.15818611337704852   0.3054019697118057   0.5671280996748016   0.18196338511525859   0.21778713677200337   0.37413422301019017   0.4834775629054257   0.06130320368273312   0.05335681452069923   0.6465784085108874   0.8565501807110518   0.5614381107757603   0.7299680258515325   0.36012588942932044   0.33824196659029376   0.6596152795812158   0.0037770635193137923   0.1906336870207076   0.7869005594999048   0.3024271197790714   0.2735759997607062   0.1308749156373558   0.7470220138927347   0.2652657094448088   0.11538988638365769   0.8254729459255501   0.17989391421793313   0.08330232432955025   0.8976027496116543   0.45133872291535987   0.6964163513125075   0.021999120646817125   0.8442459350909551   0.8047603144044724   0.8398661706014556   0.4605610098710568   0.11427790923942256   0.44463442497515193   0.5016242040111619
0.8009457302898411   0.11050084572010878   0.2540007379544444   0.7147236445112571   0.4985186105107696   0.8369248459594025   0.12312582231708857   0.9677016306185223   0.2332529010659608   0.7215349595757449   0.29765287639153853   0.7878077164005892   0.14995057673641055   0.8239322099640906   0.8463141534761787   0.09139136508808178   0.12795145608959343   0.9796862748731355   0.041553839071706226   0.25152519448662614   0.6673904462185366   0.8654083656337129   0.5969194140965542   0.7499009904754642   0.8664447159286955   0.7549075199136042   0.3429186761421099   0.03517734596420718   0.367926105417926   0.9179826739542015   0.21979285382502134   0.06747571534568483   0.13467320435196514   0.19644771437845668   0.9221399774334829   0.27966799894509564   0.9847226276155546   0.3725155044143661   0.07582582395730417   0.18827663385701385   0.8567711715259612   0.3928292295412306   0.03427198488559794   0.9367514393703876   0.18938072530742456   0.5274208639075177   0.43735257078904366   0.18685044889492342   0.32293600937872896   0.7725133439939136   0.09443389464693376   0.15167310293071623   0.955009903960803   0.854530670039712   0.8746410408219124   0.08419738758503141   0.8203366996088378   0.6580829556612553   0.9525010633884297   0.8045293886399358   0.8356140719932833   0.2855674512468892   0.8766752394311255   0.616252754782922
0.9788429004673221   0.8927382217056585   0.8424032545455274   0.6795013154125343   0.7894621751598976   0.3653173577981409   0.40505068375648384   0.49265086651761086   0.46652616578116857   0.5928040138042273   0.31061678910955004   0.34097776358689463   0.5115162618203656   0.7382733437645154   0.43597574828763763   0.2567803760018632   0.6911795622115277   0.08019038810326004   0.48347468489920803   0.4522509873619274   0.8555654902182445   0.7946229368563709   0.6067994454680826   0.8359982325790054   0.8767225897509223   0.9018847151507122   0.7643961909225551   0.15649691716647116   0.08726041459102479   0.5365673573525714   0.3593455071660713   0.6638460506488603   0.6207342488098562   0.943763343548344   0.048728718056521195   0.3228682870619657   0.10921798698949066   0.2054899997838287   0.6127529697688836   0.06608791106010248   0.418038424777963   0.12529961168056866   0.12927828486967552   0.6138369236981751   0.5624729345597186   0.3306766748241978   0.5224788394015929   0.7778386911191696   0.6857503448087962   0.42879195967348555   0.7580826484790378   0.6213417739526984   0.5984899302177714   0.8922246023209142   0.39873714131296656   0.9574957233038381   0.9777556814079151   0.9484612587725701   0.3500084232564454   0.6346274362418725   0.8685376944184245   0.7429712589887414   0.7372554534875618   0.56853952518177
0.45049926964046155   0.6176716473081727   0.6079771686178863   0.954702601483595   0.888026335080743   0.28699497248397493   0.08549832921629336   0.1768639103644253   0.20227599027194682   0.8582030128104894   0.3274156807372555   0.5555221364117269   0.6037860600541755   0.9659784104895752   0.9286785394242889   0.5980264131078887   0.6260303786462602   0.01751715171700505   0.5786701161678436   0.9633989768660163   0.7574926842278358   0.27454589272826363   0.8414146626802818   0.39485945168424624   0.3069934145873742   0.6568742454200909   0.23343749406239547   0.4401568502006513   0.4189670795066312   0.369879272936116   0.14793916484610212   0.263292939836226   0.2166910892346844   0.5116762601256266   0.8205234841088466   0.7077708034244992   0.6129050291805089   0.5456978496360515   0.8918449446845577   0.10974439031661042   0.9868746505342487   0.5281806979190464   0.3131748285167141   0.14634541345059418   0.22938196630641297   0.2536348051907828   0.4717601658364323   0.751485961766348   0.9223885517190388   0.5967605597706919   0.23832267177403682   0.31132911156569665   0.5034214722124075   0.2268812868345759   0.09038350692793472   0.04803617172947069   0.2867303829777232   0.7152050267089493   0.2698600228190881   0.34026536830497156   0.6738253537972142   0.16950717707289772   0.3780150781345305   0.23052097798836116
0.6869507032629656   0.6413264791538513   0.06484024961781644   0.08417556453776696   0.4575687369565526   0.3876916739630685   0.5930800837813841   0.332689602771419   0.5351801852375139   0.7909311141923766   0.35475741200734734   0.021360491205722344   0.03175871302510626   0.5640498273578007   0.2643739050794126   0.9733243194762516   0.7450283300473831   0.8488448006488515   0.9945138822603244   0.6330589511712801   0.07120297625016882   0.6793376235759537   0.6164988041257939   0.40253797318291895   0.38425227298720327   0.038011144422102475   0.5516585545079775   0.318362408645152   0.9266835360306507   0.6503194704590339   0.9585784707265934   0.985672805873733   0.39150335079313686   0.8593883562666573   0.6038210587192461   0.9643123146680106   0.3597446377680306   0.29533852890885665   0.33944715363983347   0.990987995191759   0.6147163077206476   0.44649372826000516   0.344933271379509   0.35792904402047887   0.5435133314704788   0.7671561046840514   0.7284344672537151   0.9553910708375599   0.15926105848327546   0.7291449602619489   0.17677591274573748   0.637028662192408   0.23257752245262475   0.07882548980291493   0.2181974420191441   0.651355856318675   0.8410741716594878   0.21943713353625754   0.614376383299898   0.6870435416506644   0.4813295338914572   0.9240986046274009   0.2749292296600645   0.6960555464589054
0.8666132261708097   0.47760487636739574   0.9299959582805555   0.3381265024384265   0.3230998947003309   0.7104487716833444   0.20156149102684046   0.3827354316008666   0.16383883621705547   0.9813038114213954   0.02478557828110297   0.7457067694084586   0.9312613137644307   0.9024783216184805   0.8065881362619589   0.09435091308978366   0.09018714210494286   0.683041188082223   0.1922117529620609   0.40730737143911927   0.6088576082134857   0.7589425834548221   0.9172825233019964   0.7112518249802139   0.742244382042676   0.28133770708742634   0.9872865650214409   0.3731253225417874   0.41914448734234505   0.5708889354040819   0.7857250739946005   0.9903898909409208   0.2553056511252896   0.5895851239826865   0.7609394957134975   0.24468312153246213   0.32404433736085886   0.687106802364206   0.9543513594515386   0.15033220844267847   0.233857195255916   0.004065614281982954   0.7621396064894777   0.7430248370035591   0.6249995870424304   0.24512303082716086   0.8448570831874813   0.03177301202334529   0.8827552049997545   0.9637853237397346   0.8575705181660404   0.6586476894815579   0.4636107176574094   0.39289638833565255   0.07184544417143995   0.6682577985406372   0.20830506653211983   0.8033112643529661   0.3109059484579425   0.42357467700817497   0.884260729171261   0.11620446198876012   0.3565545890064039   0.2732424685654965
0.650403533915345   0.11213884770677718   0.5944149825169263   0.5302176315619374   0.025403946872914564   0.8670158168796163   0.7495578993294449   0.49844461953859204   0.14264874187316012   0.9032304931398818   0.8919873811634045   0.8397969300570342   0.6790380242157508   0.5103341048042292   0.8201419369919646   0.171539131516397   0.47073295768363094   0.7070228404512632   0.5092359885340221   0.747964454508222   0.5864722285123699   0.5908183784625031   0.15268139952761817   0.4747219859427255   0.936068694597025   0.47867953075572583   0.5582664170106919   0.9445043543807882   0.9106647477241104   0.6116637138761095   0.8087085176812471   0.4460597348421962   0.7680160058509503   0.7084332207362277   0.9167211365178425   0.606262804785162   0.08897798163519956   0.19809911593199853   0.09657919952587794   0.43472367326876504   0.6182450239515687   0.4910762754807354   0.5873432109918558   0.686759218760543   0.031772795439198705   0.9002578970182323   0.4346618114642377   0.21203723281781753   0.0957041008421737   0.42157836626250655   0.8763953944535458   0.26753287843702933   0.18503935311806327   0.809914652386397   0.0676868767722987   0.8214731435948331   0.417023347267113   0.10148143165016926   0.1509657402544562   0.21521033880967114   0.32804536563191344   0.9033823157181707   0.05438654072857824   0.7804866655409061
0.7098003416803448   0.41230604023743533   0.46704332973672236   0.09372744678036306   0.678027546241146   0.512048143219203   0.03238151827248468   0.8816902139625455   0.5823234453989724   0.09046977695669643   0.15598612381893892   0.6141573355255162   0.39728409228090905   0.2805551245702994   0.08829924704664023   0.7926841919306831   0.9802607450137961   0.17907369292013017   0.9373335067921841   0.5774738531210118   0.6522153793818827   0.27569137720195946   0.8829469660636058   0.7969871875801058   0.9424150377015379   0.8633853369645241   0.41590363632688343   0.7032597407997427   0.26438749146039187   0.35133719374532113   0.38352211805439873   0.8215695268371972   0.6820640460614195   0.2608674167886247   0.2275359942354598   0.207412191311681   0.2847799537805104   0.9803122922183253   0.13923674718881957   0.41472799938099797   0.30451920876671434   0.8012385992981951   0.20190324039663554   0.8372541462599861   0.6523038293848317   0.5255472220962357   0.31895627433302975   0.04026695867988027   0.7098887916832938   0.6621618851317116   0.9030526380061463   0.33700721788013754   0.44550130022290185   0.31082469138639046   0.5195305199517476   0.5154376910429403   0.7634372541614823   0.04995727459776573   0.2919945257162878   0.3080254997312593   0.478657300380972   0.06964498237944046   0.15275777852746825   0.8932975003502613
0.17413809161425764   0.26840638308124537   0.9508545381308326   0.05604335409027526   0.521834262229426   0.7428591609850097   0.6318982637978029   0.015776395410394994   0.8119454705461323   0.0806972758532981   0.7288456257916566   0.6787691775302575   0.3664441703232304   0.7698725844669077   0.20931510583990898   0.16333148648731716   0.6030069161617481   0.719915309869142   0.9173205801236212   0.8553059867560578   0.12434961578077607   0.6502703274897015   0.7645628015961529   0.9620084864057965   0.9502115241665184   0.3818639444084561   0.8137082634653202   0.9059651323155212   0.4283772619370924   0.6390047834234465   0.18180999966751726   0.8901887369051262   0.6164317913909602   0.5583075075701484   0.4529643738758607   0.21141955937486878   0.2499876210677297   0.7884349231032407   0.2436492680359517   0.048088072887551625   0.6469807049059817   0.06851961323409875   0.32632868791233055   0.19278208613149378   0.5226310891252056   0.4182492857443973   0.5617658863161776   0.23077359972569725   0.5724195649586872   0.03638534133594113   0.7480576228508574   0.324808467410176   0.1440423030215948   0.39738055791249466   0.5662476231833402   0.43461973050504976   0.5276105116306347   0.8390730503423464   0.11328324930747952   0.22320017113018095   0.27762289056290496   0.05063812723910562   0.8696339812715278   0.17511209824262933
0.6306421856569233   0.9821185140050068   0.5433052933591973   0.9823300121111356   0.10801109653171764   0.5638692282606096   0.9815394070430196   0.7515564123854382   0.5355915315730304   0.5274838869246685   0.23348178419216217   0.4267479449752623   0.39154922855143565   0.1301033290121738   0.6672341610088219   0.9921282144702126   0.8639387169208009   0.2910302786698275   0.5539509117013425   0.7689280433400316   0.586315826357896   0.24039215143072187   0.6843169304298147   0.5938159450974022   0.9556736407009727   0.258273637425715   0.14101163707061737   0.6114859329862667   0.8476625441692551   0.6944044091651054   0.15947223002759775   0.8599295206008284   0.31207101259622466   0.16692052224043694   0.9259904458354355   0.43318157562556614   0.920521784044789   0.036817193228263136   0.2587562848266136   0.4410533611553536   0.05658306712398804   0.7457869145584356   0.7048053731252711   0.672125317815322   0.470267240766092   0.5053947631277138   0.020488442695456507   0.07830937271791973   0.5145936000651192   0.2471211257019988   0.8794768056248391   0.466823439731653   0.6669310558958641   0.5527167165368934   0.7200045755972414   0.6068939191308246   0.3548600432996395   0.38579619429645645   0.7940141297618057   0.17371234350525847   0.4343382592548504   0.3489790010681933   0.5352578449351921   0.7326589823499049
0.3777551921308624   0.6031920865097576   0.830452471809921   0.06053366453458289   0.9074879513647703   0.09779732338204389   0.8099640291144645   0.9822242918166632   0.3928943512996511   0.8506761976800451   0.9304872234896254   0.5154008520850102   0.725963295403787   0.29795948114315174   0.210482647892384   0.9085069329541855   0.3711032521041475   0.9121632868466952   0.4164685181305782   0.7347945894489271   0.936764992849297   0.563184285778502   0.881210673195386   0.0021356070990221805   0.5590098007184346   0.9599921992687444   0.05075820138546507   0.9416019425644393   0.6515218493536643   0.8621948758867004   0.24079417227100058   0.9593776507477761   0.25862749805401314   0.011518678206655322   0.3103069487813752   0.44397679866276596   0.5326642026502262   0.7135591970635036   0.09982430088899119   0.5354698657085805   0.16156095054607866   0.8013959102168083   0.6833557827584129   0.8006752762596534   0.2247959576967816   0.23821162443830635   0.8021451095630269   0.7985396691606311   0.665786156978347   0.27821942516956205   0.7513869081775618   0.8569377265961919   0.014264307624682672   0.4160245492828616   0.5105927359065613   0.8975600758484158   0.7556368095706696   0.4045058710762063   0.20028578712518605   0.4535832771856498   0.22297260692044338   0.6909466740127027   0.10046148623619484   0.9181134114770694
0.06141165637436473   0.8895507637958944   0.41710570347778186   0.11743813521741601   0.8366156986775831   0.651339139357588   0.614960593914755   0.31889846605678485   0.1708295416992362   0.373119714188026   0.8635736857371932   0.46196073946059296   0.15656523407455353   0.9570951649051644   0.35298094983063194   0.5644006636121771   0.400928424503884   0.552589293828958   0.15269516270544592   0.11081738642652736   0.17795581758344062   0.8616426198162555   0.05223367646925107   0.19270397494945798   0.11654416120907589   0.9720918560203611   0.6351279729914692   0.07526583973204197   0.2799284625314927   0.320752716662773   0.020167379076714186   0.7563673736752571   0.10909892083225656   0.947633002474747   0.156593693339521   0.2944066342146642   0.952533686757703   0.9905378375695826   0.803612743508889   0.7300059706024871   0.551605262253819   0.43794854374062453   0.6509175808034431   0.6191885841759597   0.3736494446703784   0.5763059239243691   0.598683904334192   0.42648460922650167   0.25710528346130257   0.6042140679040081   0.9635559313427229   0.3512187694944597   0.9771768209298098   0.28346135124123506   0.9433885522660087   0.5948513958192025   0.8680779000975533   0.33582834876648804   0.7867948589264877   0.30044476160453837   0.9155442133398501   0.34529051119690546   0.9831821154175987   0.5704387910020513
0.36393895108603114   0.9073419674562809   0.3322645346141555   0.9512502068260916   0.9902895064156527   0.3310360435319118   0.7335806302799635   0.52476559759959   0.7331842229543502   0.7268219756279037   0.7700246989372406   0.17354682810513028   0.7560074020245404   0.4433606243866686   0.8266361466712319   0.5786954322859277   0.8879295019269872   0.10753227562018058   0.03984128774474415   0.27825067068138937   0.972385288587137   0.7622417644232752   0.056659172327145506   0.707811879679338   0.6084463375011058   0.8548997969669943   0.72439463771299   0.7565616728532464   0.618156831085453   0.5238637534350824   0.9908140074330266   0.23179607525365634   0.8849726081311029   0.7970417778071787   0.220789308495786   0.05824924714852604   0.12896520610656254   0.35368115342051004   0.3941531618245542   0.47955381486259835   0.24103570417957537   0.24614887780032946   0.35431187407981   0.20130314418120898   0.2686504155924384   0.48390711337705433   0.2976527017526645   0.493491264501871   0.6602040780913326   0.6290073164100601   0.5732580640396745   0.7369295916486246   0.042047247005879494   0.10514356297497769   0.5824440566066479   0.5051335163949683   0.15707463887477657   0.308101785167799   0.3616547481108619   0.44688426924644226   0.028109432768214024   0.954420631747289   0.9675015862863078   0.9673304543838439
0.7870737285886387   0.7082717539469595   0.6131897122064978   0.7660273102026349   0.5184233129962003   0.22436464056990513   0.31553701045383326   0.272536045700764   0.8582192349048676   0.595357324159845   0.7422789464141588   0.5356064540521394   0.8161719878989881   0.49021376118486737   0.15983488980751082   0.030472937657171073   0.6590973490242116   0.18211197601706836   0.7981801416966489   0.5835886684107289   0.6309879162559976   0.2276913442697794   0.8306785554103412   0.6162582140268849   0.8439141876673589   0.5194195903228199   0.21748884320384337   0.8502309038242499   0.32549087467115867   0.2950549497529148   0.9019518327500101   0.577694858123486   0.46727163976629105   0.6996976255930698   0.15967288633585136   0.04208840407134658   0.6510996518673029   0.20948386440820244   0.9998379965283405   0.011615466414175506   0.9920023028430913   0.027371888391134084   0.20165785483169163   0.4280267980034467   0.3610143865870938   0.7996805441213547   0.3709792994213505   0.8117685839765618   0.5171001989197349   0.2802609537985347   0.15349045621750712   0.9615376801523119   0.1916093242485762   0.9852060040456199   0.251538623467497   0.3838428220288259   0.7243376844822852   0.2855083784525501   0.09186573713164564   0.34175441795747935   0.07323803261498223   0.07602451404434768   0.0920277406033051   0.3301389515433038
0.08123572977189088   0.04865262565321359   0.8903698857716135   0.9021121535398572   0.7202213431847971   0.24897208153185893   0.5193905863502629   0.09034356956329535   0.2031211442650622   0.9687111277333242   0.36590013013275585   0.1288058894109835   0.011511820016485996   0.9835051236877043   0.11436150666525886   0.7449630673821576   0.28717413553420085   0.6979967452351542   0.022495769533613222   0.40320864942467827   0.2139361029192186   0.6219722311908065   0.9304680289303081   0.07306969788137443   0.13270037314732774   0.573319605537593   0.04009814315869465   0.1709575443415173   0.41247902996253066   0.324347524005734   0.5207075568084317   0.08061397477822194   0.20935788569746847   0.3556363962724098   0.15480742667567582   0.9518080853672385   0.19784606568098245   0.37213127258470546   0.04044592001041697   0.20684501798508084   0.9106719301467816   0.6741345273495513   0.017950150476803744   0.8036363685604025   0.696735827227563   0.05216229615874476   0.08748212154649562   0.7305666706790281   0.5640354540802353   0.4788426906211518   0.04738397838780097   0.5596091263375108   0.1515564241177046   0.15449516661541782   0.5266764215793693   0.4789951515592889   0.9421985384202362   0.798858770343008   0.37186899490369346   0.5271870661920505   0.7443524727392536   0.42672749775830254   0.3314230748932765   0.32034204820696965
0.833680542592472   0.7525929704087513   0.31347292441647273   0.5167056796465671   0.13694471536490907   0.7004306742500065   0.22599080286997714   0.7861390089675389   0.5729092612846738   0.2215879836288547   0.17860682448217616   0.22652988263002805   0.42135283716696925   0.06709281701343688   0.6519304029028069   0.7475347310707391   0.4791542987467331   0.2682340466704288   0.2800614079991134   0.22034766487868865   0.7348018260074795   0.8415065489121263   0.9486383331058369   0.900005616671719   0.9011212834150073   0.08891357850337497   0.6351654086893641   0.38329993702515197   0.7641765680500983   0.38848290425336846   0.409174605819387   0.597160928057613   0.19126730676542442   0.16689492062451375   0.23056778133721087   0.370631045427585   0.7699144695984552   0.09980210361107689   0.578637378434404   0.6230963143568459   0.2907601708517221   0.8315680569406481   0.2985759704352906   0.40274864947815725   0.5559583448442427   0.9900615080285218   0.3499376373294537   0.5027430328064383   0.6548370614292354   0.9011479295251468   0.7147722286400895   0.1194430957812863   0.8906604933791371   0.5126650252717784   0.3055976228207025   0.5222821677236733   0.6993931866137126   0.3457701046472646   0.07502984148349166   0.15165112229608826   0.9294787170152575   0.2459680010361877   0.4963924630490877   0.5285548079392424
0.6387185461635354   0.41439994409553965   0.19781649261379708   0.12580615846108512   0.08276020131929271   0.4243384360670179   0.8478788552843434   0.6230631256546468   0.42792313989005737   0.523190506541871   0.13310662664425382   0.5036200298733605   0.5372626465109203   0.01052548127009273   0.8275090038235513   0.9813378621496873   0.8378694598972076   0.6647553766228281   0.7524791623400596   0.8296867398535991   0.9083907428819501   0.4187873755866404   0.256086699290972   0.30113193191435667   0.2696721967184147   0.004387431491100752   0.058270206677174904   0.17532577345327155   0.18691199539912198   0.5800489954240828   0.21039135139283152   0.5522626477986247   0.7589888555090646   0.05685848888221179   0.07728472474857769   0.04864261792526412   0.22172620899814435   0.04633300761211906   0.24977572092502637   0.0673047557755768   0.38385674910093676   0.38157763098929093   0.49729655858496674   0.23761801592197776   0.47546600621898666   0.9627902554026505   0.24120985929399474   0.9364860840076211   0.205793809500572   0.9584028239115497   0.18293965261681985   0.7611603105543495   0.01888181410145002   0.3783538284874669   0.9725483012239883   0.20889766275572483   0.2598929585923854   0.3214953396052551   0.8952635764754107   0.1602550448304607   0.03816674959424107   0.27516233199313606   0.6454878555503842   0.09295028905488391
0.6543100004933043   0.8935847010038451   0.14819129696541752   0.8553322731329062   0.17884399427431763   0.9307944456011946   0.9069814376714228   0.918846189125285   0.9730501847737456   0.9723916216896449   0.7240417850546029   0.15768587857093555   0.9541683706722957   0.594037793202178   0.7514934838306147   0.9487882158152107   0.6942754120799102   0.27254245359692286   0.856229907355204   0.78853317098475   0.6561086624856691   0.9973801216037869   0.21074205180481972   0.6955828819298661   0.0017986619923648294   0.10379542059994169   0.06255075483940217   0.8402506087969599   0.8229546677180472   0.17300097499874711   0.1555693171679794   0.9214044196716749   0.8499044829443015   0.20060935330910226   0.43152753211337647   0.7637185411007393   0.8957361122720059   0.6065715601069244   0.6800340482827618   0.8149303252855286   0.20146070019209572   0.33402910651000145   0.8238041409275578   0.02639715430077863   0.5453520377064266   0.33664898490621464   0.6130620891227382   0.33081427237091254   0.5435533757140618   0.23285356430627296   0.550511334283336   0.49056366357395265   0.7205987079960146   0.059852589307525864   0.3949420171153566   0.5691592439022778   0.870694225051713   0.8592432359984236   0.9634144850019801   0.8054407028015385   0.9749581127797071   0.2526716758914993   0.2833804367192183   0.9905103775160099
0.7734974125876113   0.9186425693814978   0.4595762957916604   0.9641132232152312   0.22814537488118475   0.5819935844752832   0.8465142066689223   0.6332989508443186   0.684591999167123   0.3491400201690102   0.2960028723855863   0.14273528727036602   0.9639932911711084   0.2892874308614843   0.9010608552702297   0.5735760433680882   0.0932990661193954   0.4300441948630607   0.9376463702682496   0.7681353405665498   0.11834095333968833   0.17737251897156142   0.6542659335490313   0.77762496305054   0.344843540752077   0.2587299495900636   0.19468963775737086   0.8135117398353087   0.11669816587089224   0.6767363651147805   0.34817543108844856   0.18021278899099005   0.4321061667037693   0.32759634494577033   0.052172558702862304   0.03747750172062401   0.46811287553266084   0.03830891408428602   0.1511117034326326   0.46390145835253577   0.3748138094132655   0.6082647192212253   0.21346533316438304   0.695766117785986   0.2564728560735771   0.4308922002496639   0.5591993996153517   0.9181411547354461   0.9116293153215002   0.17216225065960028   0.3645097618579809   0.10462941490013734   0.7949311494506079   0.4954258855448198   0.016334330769532304   0.9244166259091473   0.3628249827468386   0.16782954059904945   0.96416177206667   0.8869391241885233   0.8947121072141778   0.12952062651476343   0.8130500686340374   0.42303766583598756
0.5198982978009123   0.5212559072935381   0.5995847354696544   0.7272715480500016   0.2634254417273352   0.09036370704387423   0.04038533585430262   0.8091303933145555   0.351796126405835   0.918201456384274   0.6758755739963217   0.7045009784144182   0.5568649769552271   0.42277557083945416   0.6595412432267894   0.7800843525052709   0.1940399942083885   0.2549460302404047   0.6953794711601194   0.8931452283167476   0.29932788699421076   0.12542540372564126   0.882329402526082   0.47010756248076   0.7794295891932984   0.6041694964321032   0.28274466705642765   0.7428360144307584   0.5160041474659632   0.513805789388229   0.24235933120212502   0.9337056211162029   0.16420802106012822   0.595604333003955   0.5664837572058032   0.22920464270178478   0.6073430441049011   0.17282876216450083   0.9069425139790138   0.44912029019651395   0.4133030498965126   0.9178827319240961   0.21156304281889443   0.5559750618797664   0.11397516290230186   0.7924573281984548   0.32923364029281244   0.0858674993990064   0.33454557370900345   0.1882878317663517   0.04648897323638477   0.3430314849682479   0.8185414262430402   0.6744820423781228   0.8041296420342597   0.409325863852045   0.6543334051829119   0.0788777093741678   0.23764588482845644   0.1801212211502602   0.04699036107801085   0.906048947209667   0.33070337084944257   0.7310009309537463
0.6336873111814982   0.9881662152855709   0.11914032803054816   0.17502586907397985   0.5197121482791964   0.195708887087116   0.7899066877377358   0.08915836967497345   0.18516657457019298   0.0074210553207643085   0.743417714501351   0.7461268847067255   0.3666251483271528   0.33293901294264155   0.9392880724670912   0.3368010208546805   0.7122917431442408   0.25406130356847373   0.7016421876386347   0.15667979970442034   0.66530138206623   0.34801235635880673   0.3709388167891922   0.42567886875067407   0.03161407088473174   0.35984614107323587   0.251798488758644   0.25065299967669424   0.5119019226055354   0.16413725398611986   0.46189180102090827   0.16149463000172076   0.3267353480353424   0.15671619866535555   0.7184740865195574   0.41536774529499526   0.9601101997081896   0.8237771857227141   0.779186014052466   0.07856672444031475   0.2478184565639487   0.5697158821542403   0.07754382641383128   0.9218869247358944   0.5825170744977187   0.22170352579543356   0.7066050096246391   0.49620805598522033   0.5509030036129869   0.8618573847221976   0.45480652086599505   0.24555505630852612   0.03900108100745166   0.6977201307360779   0.9929147198450868   0.08406042630680534   0.7122657329721093   0.5410039320707223   0.2744406333255295   0.6686926810118101   0.7521555332639197   0.7172267463480082   0.4952546192730634   0.5901259565714954
0.504337076699971   0.14751086419376794   0.4177107928592321   0.668239031835601   0.9218200022022522   0.9258073383983344   0.7111057832345931   0.17203097585038057   0.37091699858926525   0.0639499536761367   0.25629926236859796   0.9264759195418545   0.3319159175818136   0.3662298229400589   0.2633845425235112   0.8424154932350492   0.6196501846097043   0.8252258908693366   0.9889439091979817   0.17372281222323904   0.8674946513457846   0.10799914452132842   0.4936892899249183   0.5835968556517437   0.3631575746458136   0.9604882803275605   0.07597849706568617   0.9153578238161428   0.44133757244356137   0.0346809419292261   0.36487271383109315   0.7433268479657622   0.07042057385429609   0.9707309882530893   0.1085734514624952   0.8168509284239077   0.7385046562724825   0.6045011653130304   0.845188908938984   0.9744354351888587   0.11885447166277817   0.7792752744436938   0.8562449997410023   0.8007126229656196   0.25135982031699355   0.6712761299223654   0.36255570981608404   0.21711576731387588   0.8882022456711799   0.7107878495948049   0.2865772127503979   0.3017579434977331   0.4468646732276186   0.6761069076655789   0.9217044989193047   0.5584310955319709   0.37644409937332246   0.7053759194124894   0.8131310474568095   0.7415801671080631   0.63793944310084   0.10087475409945897   0.9679421385178255   0.7671447319192045
0.5190849714380619   0.32159947965576513   0.11169713877682319   0.9664321089535849   0.26772515112106826   0.6503233497333997   0.7491414289607392   0.749316341639709   0.3795229054498883   0.9395355001385948   0.46256421621034133   0.4475583981419759   0.9326582322222697   0.26342859247301587   0.5408597172910365   0.889127302610005   0.5562141328489473   0.5580526730605264   0.7277286698342271   0.1475471355019419   0.9182746897481072   0.45717791896106746   0.7597865313164016   0.3804024035827374   0.39918971831004546   0.13557843930530233   0.6480893925395784   0.4139702946291525   0.13146456718897717   0.48525508957190266   0.8989479635788392   0.6646539529894435   0.7519416617390888   0.5457195894333079   0.43638374736849794   0.21709555484746765   0.8192834295168191   0.2822909969602921   0.8955240300774613   0.3279682522374626   0.2630692966678718   0.7242383238997656   0.16779536024323424   0.18042111673552072   0.34479460691976455   0.2670604049386982   0.40800882892683266   0.8000187131527833   0.9456048886097191   0.13148196563339587   0.7599194363872542   0.3860484185236307   0.8141403214207419   0.6462268760614932   0.860971472808415   0.7213944655341872   0.062198659681653105   0.10050728662818527   0.42458772543991713   0.5042989106867195   0.24291523016483405   0.8182162896678932   0.5290636953624558   0.17633065844925688
0.9798459334969623   0.09397796576812754   0.3612683351192216   0.9959095417137361   0.6350513265771978   0.8269175608294294   0.9532595061923889   0.1958908285609529   0.6894464379674786   0.6954355951960335   0.19334006980513457   0.8098424100373222   0.8753061165467367   0.049208719134540245   0.33236859699671956   0.088447944503135   0.8131074568650836   0.948701432506355   0.9077808715568024   0.5841490338164155   0.5701922267002495   0.13048514283846177   0.3787171761943466   0.4078183753671586   0.5903462932032874   0.03650717707033425   0.017448841075125055   0.4119088336534224   0.9552949666260896   0.2095896162409049   0.06418933488273618   0.2160180050924695   0.26584852865861097   0.5141540210448715   0.8708492650776016   0.40617559505514733   0.39054241211187424   0.46494530191033123   0.538480668080882   0.3177276505520123   0.5774349552467907   0.5162438694039763   0.6306997965240797   0.7335786167355968   0.00724272854654112   0.38575872656551446   0.25198262032973306   0.32576024136843823   0.4168964353432538   0.3492515494951802   0.234533779254608   0.9138514077150158   0.46160146871716423   0.13966193325427528   0.17034444437187182   0.6978334026225463   0.1957529400585533   0.6255079122094038   0.2994951792942702   0.291657807567399   0.805210527946679   0.16056261029907262   0.7610145112133881   0.9739301570153867
0.22777557269988835   0.6443187408950964   0.1303147146893085   0.24035154027978986   0.22053284415334723   0.2585600143295819   0.8783320943595755   0.9145912989113516   0.8036364088100935   0.9093084648344018   0.6437983151049674   0.000739891196335845   0.3420349400929292   0.7696465315801264   0.47345387073309564   0.30290648857378955   0.14628200003437591   0.14413861937072261   0.1739586914388254   0.011248681006390558   0.3410714720876969   0.98357600907165   0.4129441802254372   0.037318523991003875   0.11329589938780854   0.3392572681765536   0.2826294655361287   0.796966983711214   0.8927630552344613   0.08069725384697167   0.4042973711765533   0.8823756847998624   0.0891266464243679   0.17138878901256993   0.7604990560715859   0.8816357936035265   0.7470917063314387   0.40174225743244346   0.28704518533849027   0.578729305029737   0.6008097062970628   0.2576036380617208   0.11308649389966485   0.5674806240233464   0.2597382342093659   0.2740276289900708   0.7001423136742276   0.5301621000323425   0.14644233482155739   0.9347703608135172   0.41751284813809886   0.7331951163211285   0.2536792795870961   0.8540731069665456   0.013215476961545566   0.8508194315212662   0.16455263316272817   0.6826843179539757   0.2527164208899597   0.9691836379177396   0.41746092683128944   0.28094206052153214   0.9656712355514695   0.3904543328880027
0.8166512205342267   0.023338422459811325   0.8525847416518046   0.8229737088646563   0.5569129863248607   0.7493107934697405   0.15244242797757698   0.2928116088323137   0.4104706515033033   0.8145404326562232   0.7349295798394782   0.5596164925111852   0.15679137191620726   0.9604673256896777   0.7217141028779326   0.708797060989919   0.9922387387534791   0.2777830077357021   0.46899768198797287   0.7396134230721794   0.5747778119221897   0.9968409472141699   0.5033264464365034   0.3491590901841767   0.758126591387963   0.9735025247543586   0.6507417047846988   0.5261853813195204   0.2012136050631023   0.2241917312846181   0.4982992768071218   0.23337377248720673   0.790742953559799   0.40965129862839483   0.7633696969676437   0.6737572799760215   0.6339515816435917   0.4491839729387171   0.04165559408971116   0.9649602189861025   0.6417128428901127   0.171400965203015   0.5726579121017383   0.22534679591392312   0.06693503096792297   0.17456001798884507   0.06933146566523492   0.8761877057297465   0.30880843957995996   0.20105749323448646   0.4185897608805361   0.350002324410226   0.10759483451685768   0.9768657619498684   0.9202904840734143   0.11662855192301926   0.31685188095705874   0.5672144633214735   0.1569207871057706   0.4428712719469977   0.6829002993134671   0.1180304903827564   0.11526519301605943   0.4779110529608952
0.04118745642335443   0.9466295251797414   0.5426072809143211   0.2525642570469721   0.9742524254554314   0.7720695071908963   0.4732758152490862   0.37637655131722564   0.6654439858754715   0.5710120139564098   0.0546860543685501   0.026374226906999674   0.5578491513586138   0.5941462520065415   0.1343955702951358   0.9097456749839804   0.2409972704015551   0.02693178868506795   0.9774747831893652   0.4668744030369827   0.5580969710880881   0.9089012983023116   0.8622095901733058   0.9889633500760875   0.5169095146647337   0.9622717731225702   0.31960230925898464   0.7363990930291154   0.5426570892093021   0.1902022659316739   0.8463264940098985   0.36002254171188974   0.8772131033338306   0.6191902519752641   0.7916404396413483   0.3336483148048901   0.31936395197521683   0.0250439999687226   0.6572448693462125   0.42390263982090964   0.07836668157366174   0.9981122112836547   0.6797700861568473   0.957028236783927   0.5202697104855737   0.0892109129813431   0.8175604959835415   0.9680648867078394   0.003360195820840052   0.12693913985877292   0.4979581867245569   0.23166579367872406   0.4607031066115379   0.936736873927099   0.6516316927146585   0.8716432519668342   0.5834900032777073   0.317546621951835   0.85999125307331   0.5379949371619442   0.2641260513024904   0.2925026219831124   0.20274638372709752   0.11409229734103453
0.18575936972882864   0.2943904106994577   0.5229762975702502   0.1570640605571076   0.665489659243255   0.20517949771811464   0.7054158015867086   0.18899917384926812   0.662129463422415   0.07824035785934172   0.20745761486215172   0.957333380170544   0.20142635681087703   0.14150348393224269   0.5558259221474933   0.08569012820370978   0.6179363535331698   0.8239568619804077   0.6958346690741832   0.5476951910417656   0.3538103022306794   0.5314542399972954   0.49308828534708565   0.4336028937007311   0.16805093250185077   0.2370638292978376   0.9701119877768355   0.2765388331436235   0.5025612732585958   0.03188433157972295   0.26469618619012686   0.08753965929435537   0.8404318098361808   0.9536439737203812   0.057238571327975156   0.1302062791238113   0.6390054530253039   0.8121404897881386   0.5014126491804819   0.04451615092010152   0.02106909949213405   0.9881836278077308   0.8055779801062987   0.4968209598783359   0.6672587972614547   0.45672938781043554   0.31248969475921307   0.06321806617760489   0.4992078647596039   0.21966555851259795   0.34237770698237757   0.7866792330339815   0.9966465915010081   0.187781226932875   0.0776815207922507   0.6991395737396261   0.15621478166482722   0.23413725321249376   0.020442949464275537   0.5689332946158148   0.5172093286395234   0.4219967634243552   0.5190303002837936   0.5244171436957132
0.4961402291473893   0.4338131356166243   0.7134523201774949   0.027596183817377298   0.8288814318859347   0.9770837478061888   0.40096262541828187   0.9643781176397724   0.3296735671263308   0.7574181892935908   0.05858491843590433   0.177698884605791   0.3330269756253227   0.5696369623607158   0.9809033976436536   0.47855931086616493   0.17681219396049547   0.3354997091482221   0.9604604481793781   0.9096260162503502   0.6596028653209721   0.9135029457238669   0.44143014789558443   0.3852088725546369   0.16346263617358275   0.47968981010724254   0.7279778277180895   0.35761268873725965   0.33458120428764804   0.5026060623010538   0.32701520229980763   0.3932345710974872   0.004907637161317272   0.7451878730074629   0.2684302838639033   0.21553568649169624   0.6718806615359946   0.17555091064674705   0.28752688622024963   0.7369763756255313   0.4950684675754991   0.840051201498525   0.32706643804087154   0.8273503593751811   0.835465602254527   0.926548255774658   0.8856362901452871   0.44214148682054416   0.6720029660809443   0.4468584456674155   0.15765846242719758   0.08452879808328453   0.33742176179329625   0.9442523833663617   0.83064326012739   0.6912942269857973   0.33251412463197894   0.19906451035889886   0.5622129762634867   0.47575854049410105   0.6606334630959844   0.02351359971215181   0.274686090043237   0.7387821648685697
0.16556499552048526   0.18346239821362684   0.9476196520023654   0.9114318054933886   0.3300993932659582   0.25691414243896876   0.06198336185707838   0.46929031867284443   0.6580964271850139   0.8100556967715532   0.9043248994298808   0.3847615205895599   0.3206746653917177   0.8658033134051915   0.07368163930249086   0.6934672936037626   0.9881605407597387   0.6667388030462926   0.5114686630390042   0.21770875310966156   0.3275270776637544   0.6432252033341408   0.2367825729957672   0.47892658824109186   0.1619620821432691   0.459762805120514   0.28916292099340174   0.5674947827477033   0.8318626888773109   0.2028486626815452   0.22717955913632334   0.09820446407485876   0.17376626169229697   0.39279296590999196   0.32285465970644256   0.7134429434852988   0.8530915963005793   0.5269896525048005   0.24917302040395167   0.01997564988153623   0.8649310555408406   0.8602508494585078   0.7377043573649474   0.8022668967718747   0.5374039778770862   0.21702564612436703   0.5009217843691803   0.3233403085307828   0.3754418957338171   0.7572628410038531   0.21175886337577857   0.7558455257830796   0.5435792068565062   0.5544141783223079   0.9845793042394552   0.6576410617082209   0.3698129451642092   0.16162121241231595   0.6617246445330127   0.944198118222922   0.51672134886363   0.6346315599075155   0.412551624129061   0.9242224683413858
0.6517902933227894   0.7743807104490076   0.6748472667641136   0.1219555715695111   0.11438631544570316   0.5573550643246405   0.17392548239493325   0.7986152630387283   0.7389444197118861   0.8000922233207876   0.9621666190191547   0.042769737255648664   0.19536521285537986   0.24567804499847962   0.9775873147796995   0.3851286755474278   0.8255522676911706   0.08405683258616366   0.3158626702466868   0.4409305573245058   0.3088309188275407   0.4494252726786482   0.9033110461176258   0.51670808898312   0.6570406255047514   0.6750445622296405   0.22846377935351228   0.39475251741360895   0.5426543100590482   0.11768949790499994   0.05453829695857903   0.5961372543748806   0.8037098903471621   0.31759727458421244   0.09237167793942434   0.553367517119232   0.6083446774917823   0.07191922958573284   0.11478436315972487   0.1682388415718042   0.7827924098006116   0.9878623969995691   0.798921692913038   0.7273082842472983   0.47396149097307094   0.5384371243209211   0.8956106467954122   0.2106001952641783   0.8169208654683195   0.8633925620912805   0.6671468674419   0.8158476778505693   0.27426655540927136   0.7457030641862805   0.612608570483321   0.2197104234756887   0.4705566650621092   0.4281057896020681   0.5202368925438966   0.6663429063564567   0.8622119875703269   0.35618656001633525   0.40545252938417176   0.4981040647846525
0.07941957776971525   0.36832416301676607   0.6065308364711337   0.7707957805373542   0.6054580867966444   0.829887038695845   0.7109201896757215   0.5601955852731758   0.7885372213283248   0.9664944766045646   0.04377332223382142   0.7443479074226065   0.5142706659190535   0.22079141241828407   0.43116475175050045   0.5246374839469178   0.04371400085694424   0.792685622816216   0.9109278592066038   0.8582945775904611   0.18150201328661733   0.4364990627998807   0.505475329822432   0.3601905128058086   0.10208243551690209   0.06817489978311465   0.8989444933512983   0.5893947322684544   0.49662434872025774   0.2382878610872696   0.1880243036755769   0.029199146995278587   0.708087127391933   0.271793384482705   0.1442509814417555   0.28485123957267205   0.19381646147287954   0.051001972064420954   0.713086229691255   0.7602137556257542   0.1501024606159353   0.258316349248205   0.8021583704846512   0.9019191780352932   0.9686004473293179   0.8218172864483243   0.29668304066221923   0.5417286652294846   0.8665180118124158   0.7536423866652097   0.3977385473109209   0.9523339329610301   0.3698936630921581   0.51535452557794   0.20971424363534397   0.9231347859657515   0.6618065357002252   0.24356114109523502   0.06546326219358849   0.6382835463930794   0.46799007422734556   0.19255916903081408   0.35237703250233343   0.8780697907673252
0.31788761361141027   0.934242819782609   0.5502186620176822   0.976150612732032   0.34928716628209233   0.11242553333428482   0.253535621355463   0.4344219475025475   0.48276915446967644   0.3587831466690752   0.8557970740445421   0.4820880145415174   0.11287549137751833   0.8434286210911351   0.6460828304091981   0.5589532285757659   0.4510689556772932   0.5998674799959002   0.5806195682156097   0.9206696821826864   0.9830788814499476   0.4073083109650861   0.22824253571327618   0.04259989141536127   0.6651912678385373   0.473065491182477   0.678023873695594   0.06644927868332925   0.315904101556445   0.3606399578481922   0.424488252340131   0.6320273311807818   0.8331349470867686   0.001856811179116976   0.5686911782955889   0.1499393166392644   0.7202594557092502   0.1584281900879818   0.9226083478863908   0.5909860880634985   0.26919050003195705   0.5585607100920816   0.3419887796707812   0.6703164058808121   0.2861116185820094   0.1512523991269956   0.113746243957505   0.6277165144654508   0.6209203507434721   0.6781869079445186   0.435722370261911   0.5612672357821216   0.3050162491870271   0.31754695009632644   0.011234117921780022   0.9292399046013398   0.4718813021002585   0.31569013891720943   0.4425429396261911   0.7793005879620754   0.7516218463910083   0.15726194882922764   0.5199345917398003   0.18831449989857685
0.4824313463590512   0.598701238737146   0.17794581206901913   0.5179980940177648   0.19631972777704182   0.44744883961015036   0.06419956811151412   0.8902815795523139   0.5753993770335697   0.7692619316656318   0.6284771978496031   0.3290143437701923   0.27038312784654267   0.45171498156930534   0.6172430799278231   0.39977443916885247   0.7985018257462841   0.1360248426520959   0.17470014030163197   0.6204738512067771   0.04687997935527588   0.9787628938228683   0.6547655485618317   0.43215935130820027   0.5644486329962246   0.38006165508572226   0.4768197364928125   0.9141612572904355   0.36812890521918284   0.9326128154755718   0.4126201683812984   0.023879677738121628   0.792729528185613   0.16335088380994012   0.7841429705316953   0.6948653339679294   0.5223464003390704   0.7116359022406348   0.16689989060387225   0.29509089479907685   0.7238445745927863   0.5756110595885389   0.9921997503022403   0.6746170435922998   0.6769645952375104   0.5968481657656706   0.3374342017404086   0.24245769228409952   0.11251596224128575   0.2167865106799483   0.8606144652475961   0.328296434993664   0.744387057022103   0.2841736952043764   0.44799429686629766   0.30441675725554235   0.9516575288364899   0.12082281139443629   0.6638513263346024   0.609551423287613   0.4293111284974194   0.4091869091538015   0.49695143573073014   0.3144605284885362
0.7054665539046332   0.8335758495652626   0.5047516854284898   0.6398434848962364   0.028501958667122754   0.2367276837995921   0.16731748368808122   0.3973857926121369   0.915985996425837   0.01994117311964381   0.30670301844048514   0.06908935761847292   0.17159893940373405   0.7357674779152674   0.8587087215741874   0.7646726003629305   0.2199414105672442   0.6149446665208311   0.19485739523958506   0.1551211770753175   0.7906302820698248   0.2057577573670296   0.6979059595088549   0.8406606485867814   0.08516372816519162   0.3721819078017669   0.1931542740803651   0.2008171636905449   0.05666176949806887   0.1354542240021748   0.02583679039228388   0.803431371078408   0.14067577307223186   0.11551305088253098   0.7191337719517987   0.734342013459935   0.9690768336684978   0.3797455729672636   0.8604250503776113   0.9696694130970045   0.7491354231012536   0.7648009064464325   0.6655676551380263   0.814548236021687   0.9585051410314288   0.5590431490794029   0.9676616956291714   0.9738875874349057   0.8733414128662372   0.18686124127763598   0.7745074215488063   0.7730704237443607   0.8166796433681683   0.05140701727546119   0.7486706311565223   0.9696390526659528   0.6760038702959364   0.9358939663929302   0.02953685920472359   0.2352970392060178   0.7069270366274386   0.5561483934256666   0.16911180882711227   0.2656276261090133
0.957791613526185   0.7913474869792342   0.503544153689086   0.4510793900873263   0.9992864724947562   0.2323043378998313   0.5358824580599146   0.4771918026524206   0.12594505962851898   0.045443096622195325   0.7613750365111084   0.7041213789080598   0.30926541626035065   0.9940360793467341   0.012704405354586064   0.734482326242107   0.6332615459644142   0.05814211295380393   0.9831675461498625   0.49918528703608916   0.9263345093369755   0.5019937195281373   0.8140557373227502   0.2335576609270759   0.9685428958107904   0.7106462325489031   0.3105115836336642   0.7824782708397496   0.9692564233160342   0.47834189464907184   0.7746291255737495   0.30528646818732896   0.8433113636875154   0.4328987980268765   0.013254089062641142   0.6011650892792691   0.5340459474271647   0.43886271868014237   0.0005496837080550773   0.8666827630371622   0.9007844014627505   0.3807206057263384   0.017382137558192606   0.36749747600107296   0.974449892125775   0.8787268861982012   0.2033264002354424   0.13393981507399708   0.00590699631498455   0.168080653649298   0.8928148166017782   0.3514615442342475   0.03665057299895027   0.6897387590002262   0.11818569102802862   0.046175076046918534   0.19333920931143495   0.2568399609733497   0.10493160196538746   0.4450099867676494   0.6592932618842703   0.8179772422932073   0.1043819182573324   0.5783272237304872
0.7585088604215198   0.4372566365668689   0.08699978069913979   0.21082974772941424   0.7840589682957447   0.5585297503686678   0.8836733804636974   0.07688993265541716   0.7781519719807601   0.3904490967193698   0.9908585638619192   0.7254283884211696   0.7415013989818099   0.7007103377191436   0.8726728728338906   0.6792533123742511   0.548162189670375   0.4438703767457939   0.7677412708685032   0.23424332560660174   0.8888689277861047   0.6258931344525865   0.6633593526111707   0.6559161018761145   0.13036006736458491   0.18863649788571765   0.5763595719120309   0.4450863541467003   0.3463010990688402   0.6301067475170499   0.6926861914483335   0.3681964214912831   0.56814912708808   0.23965765079768012   0.7018276275864144   0.6427680330701134   0.8266477281062701   0.5389473130785365   0.8291547547525238   0.9635147206958623   0.27848553843589513   0.09507693633274265   0.061413483884020605   0.7292713950892605   0.3896166106497905   0.46918380188015607   0.39805413127284983   0.07335529321314607   0.25925654328520553   0.28054730399443845   0.8216945593608189   0.6282689390664458   0.9129554442163653   0.6504405564773885   0.12900836791248532   0.2600725175751627   0.34480631712828536   0.41078290567970843   0.42718074032607095   0.6173044845050493   0.5181585890220153   0.8718355926011718   0.5980259855735472   0.653789763809187
0.23967305058612007   0.7767586562684292   0.5366125016895267   0.9245183687199263   0.8500564399363296   0.30757485438827314   0.13855837041667676   0.8511630755067803   0.5907998966511241   0.027027550393834712   0.31686381105585787   0.22289413644033448   0.6778444524347587   0.3765869939164462   0.18785544314337255   0.9628216188651718   0.3330381353064733   0.9658040882367378   0.7606747028173015   0.34551713436012255   0.8148795462844581   0.09396849563556592   0.16264871724375435   0.6917273705509356   0.575206495698338   0.3172098393671367   0.6260362155542277   0.7672090018310093   0.7251500557620084   0.009634984978863562   0.48747784513755094   0.916045926324229   0.13435015911088438   0.9826074345850289   0.17061403408169307   0.6931517898838945   0.4565057066761257   0.6060204406685826   0.9827585909383205   0.7303301710187227   0.12346757136965239   0.6402163524318449   0.22208388812101898   0.38481303665860017   0.3085880250851943   0.546247856796279   0.059435170877264645   0.6930856661076645   0.7333815293868563   0.2290380174291423   0.4333989553230369   0.9258766642766554   0.008231473624847859   0.21940303245027873   0.945921110185486   0.009830737952426396   0.8738813145139634   0.23679559786524987   0.7753070761037929   0.3166789480685319   0.4173756078378378   0.6307751571966672   0.7925484851654724   0.5863487770498093
0.29390803646818536   0.9905588047648223   0.5704645970444534   0.20153574039120906   0.9853200113829911   0.44431094796854337   0.5110294261671887   0.5084500742835445   0.25193848199613483   0.21527293053940105   0.07763047084415181   0.5825734100068891   0.24370700837128695   0.9958698980891223   0.13170936065866581   0.5727426720544627   0.36982569385732345   0.7590743002238725   0.35640228455487294   0.2560637239859308   0.9524500860194857   0.12829914302720527   0.5638537993894006   0.6697149469361215   0.6585420495513004   0.13774033826238297   0.9933892023449472   0.4681792065449125   0.6732220381683093   0.6934293902938397   0.48235977617775844   0.959729132261368   0.42128355617217444   0.47815645975443855   0.4047293053336066   0.3771557222544789   0.1775765478008875   0.4822865616653162   0.2730199446749408   0.8044130502000162   0.807750853943564   0.7232122614414437   0.9166176601200678   0.5483493262140854   0.8553007679240783   0.5949131184142384   0.3527638607306673   0.8786343792779638   0.19675871837277797   0.4571727801518555   0.35937465838572014   0.41045517273305127   0.5235366802044688   0.7637433898580158   0.8770148822079618   0.45072604047168324   0.10225312403229429   0.2855869301035773   0.4722855768743551   0.07357031821720429   0.9246765762314068   0.8033003684382611   0.1992656321994143   0.2691572680171881
0.11692572228784279   0.08008810699681737   0.28264797207934644   0.7208079418031027   0.2616249543637645   0.48517498858257896   0.9298841113486791   0.842173562525139   0.0648662359909865   0.028002208430723464   0.570509452962959   0.43171838979208765   0.5413295557865178   0.2642588185727076   0.6934945707549972   0.9809923493204045   0.43907643175422345   0.9786718884691303   0.22120899388064216   0.9074220311032002   0.5143998555228166   0.17537152003086923   0.021943361681227885   0.6382647630860121   0.3974741332349739   0.09528341303405184   0.7392953896018815   0.9174568212829093   0.1358491788712094   0.610108424451473   0.8094112782532024   0.07528325875777037   0.07098294288022292   0.5821062160207494   0.2389018252902434   0.6435648689656827   0.5296533870937051   0.3178473974480418   0.5454072545352462   0.6625725196452782   0.09057695533948168   0.3391755089789115   0.32419826065460394   0.7551504885420781   0.576177099816665   0.1638039889480423   0.3022548989733761   0.116885725456066   0.17870296658169113   0.06852057591399047   0.5629595093714946   0.1994289041731567   0.04285378771048172   0.45841215146251757   0.7535482311182923   0.12414564541538632   0.9718708448302588   0.8763059354417682   0.5146464058280489   0.48058077644970365   0.44221745773655363   0.5584585379937264   0.9692391512928027   0.8180082568044253
0.35164050239707195   0.21928302901481478   0.6450408906381988   0.06285776826234733   0.7754634025804069   0.05547904006677249   0.3427859916648227   0.9459720428062813   0.5967604359987159   0.986958464152782   0.7798264822933281   0.7465431386331246   0.5539066482882341   0.5285463126902644   0.02627825117503583   0.6223974932177383   0.5820358034579753   0.6522403772484964   0.511631845346987   0.1418167167680347   0.13981834572142166   0.09378183925477002   0.5423926940541842   0.3238084599636093   0.7881778433243497   0.8744988102399552   0.8973518034159855   0.26095069170126195   0.012714440743942712   0.8190197701731827   0.5545658117511628   0.3149786488949806   0.41595400474522687   0.8320613060204007   0.7747393294578347   0.568435510261856   0.8620473564569928   0.30351499333013626   0.748461078282799   0.9460380170441176   0.2800115529990175   0.65127461608164   0.23682923293581193   0.804221300276083   0.14019320727759582   0.5574927768268699   0.6944365388816277   0.48041284031247367   0.3520153639532461   0.6829939665869147   0.7970847354656422   0.2194621486112117   0.33930092320930344   0.863974196413732   0.24251892371447936   0.9044834997162311   0.9233469184640766   0.03191289039333124   0.46777959425664467   0.3360479894543751   0.06129956200708378   0.728397897063195   0.7193185159738458   0.3900099724102574
0.7812880090080663   0.07712328098155503   0.48248928303803384   0.5857886721341745   0.6410948017304705   0.5196305041546851   0.7880527441564061   0.10537583182170081   0.2890794377772244   0.8366365375677705   0.990968008690764   0.8859136832104891   0.949778514567921   0.9726623411540385   0.7484490849762846   0.981430183494258   0.026431596103844386   0.9407494507607073   0.2806694907196399   0.645382194039883   0.9651320340967606   0.21235155369751224   0.5613509747457942   0.25537222162962553   0.1838440250886943   0.1352282727159572   0.07886169170776038   0.6695835494954511   0.5427492233582237   0.6155977685612721   0.2908089475513542   0.5642077176737503   0.2536697855809994   0.7789612309935017   0.29984093886059027   0.6782940344632612   0.3038912710130785   0.8062988898394632   0.5513918538843057   0.6968638509690032   0.27745967490923407   0.865549439078756   0.27072236316466575   0.05148165692912016   0.3123276408124735   0.6531978853812438   0.7093713884188716   0.7961094352994946   0.1284836157237792   0.5179696126652865   0.6305096967111111   0.12652588580404353   0.5857343923655555   0.9023718441040145   0.33970074915975695   0.5623181681302932   0.332064606784556   0.12341061311051278   0.039859810299166666   0.8840241336670321   0.02817333577147754   0.3171117232710496   0.48846795641486096   0.18716028269802898
0.7507136608622434   0.4515622841922936   0.21774559325019524   0.13567862576890882   0.43838602004976995   0.7983643988110498   0.5083742048313237   0.3395691904694142   0.30990240432599075   0.2803947861457633   0.8778645081202125   0.21304330466537064   0.7241680119604353   0.3780229420417488   0.5381637589604555   0.6507251365350774   0.39210340517587927   0.25461232893123603   0.4983039486612889   0.7667010028680453   0.36393006940440176   0.9375006056601864   0.00983599224642793   0.5795407201700163   0.6132164085421583   0.4859383214678929   0.7920903989962327   0.4438620944011075   0.17483038849238836   0.687573922656843   0.283716194164909   0.10429290393169331   0.8649279841663976   0.4071791365110798   0.40585168604469646   0.8912495992663226   0.14075997220596229   0.029156194469330942   0.8676879270842409   0.24052446273124528   0.748656567030083   0.774543865538095   0.36938397842295195   0.4738234598632   0.38472649762568123   0.8370432598779085   0.35954798617652406   0.8942827396931837   0.7715100890835229   0.35110493841001555   0.5674575871802914   0.4504206452920762   0.5966797005911346   0.6635310157531725   0.28374139301538237   0.3461277413603829   0.731751716424737   0.2563518792420928   0.8778897069706859   0.4548781420940602   0.5909917442187747   0.22719568477276184   0.010201779886445009   0.21435367936281494
0.8423351771886917   0.4526518192346669   0.6408178014634931   0.740530219499615   0.45760867956301043   0.6156085593567585   0.281269815286969   0.8462474798064312   0.6860985904794875   0.2645036209467429   0.7138122281066777   0.3958268345143551   0.08941888988835292   0.6009726051935703   0.4300708350912953   0.04969909315397223   0.357667173463616   0.3446207259514776   0.5521811281206094   0.5948209510599121   0.7666754292448413   0.11742504117871576   0.5419793482341644   0.3804672716970971   0.9243402520561497   0.6647732219440489   0.9011615467706714   0.6399370521974821   0.4667315724931392   0.049164662587290374   0.6198917314837024   0.7936895723910509   0.7806329820136517   0.7846610416405475   0.9060795033770247   0.39786273787669574   0.6912140921252987   0.18368843644697713   0.4760086682857294   0.3481636447227235   0.3335469186616828   0.8390677104954996   0.92382754016512   0.7533426936628115   0.5668714894168415   0.7216426693167838   0.3818481919309556   0.37287542196571444   0.6425312373606918   0.056869447372734944   0.4806866451602842   0.7329383697682323   0.1757996648675527   0.0077047847854445715   0.8607949136765819   0.9392487973771815   0.395166682853901   0.22304374314489708   0.9547154102995572   0.5413860595004857   0.7039525907286023   0.03935530669791995   0.4787067420138278   0.19322241477776222
0.37040567206691943   0.2002875962024204   0.5548792018487079   0.4398797211149507   0.8035341826500779   0.47864492688563665   0.17303100991775225   0.0670042991492363   0.16100294528938605   0.4217754795129017   0.6923443647574681   0.334065929381004   0.9852032804218334   0.4140706947274571   0.8315494510808862   0.3948171320038225   0.5900365975679324   0.19102695158256003   0.876834040781329   0.8534310725033368   0.8860840068393301   0.15167164488464008   0.3981272987675012   0.6602086577255746   0.5156783347724107   0.9513840486822197   0.8432480969187933   0.22032893661062386   0.7121441521223327   0.472739121796583   0.6702170870010411   0.15332463746138758   0.5511412068329467   0.05096364228368136   0.9778727222435731   0.8192587080803836   0.5659379264111133   0.6368929475562243   0.14632327116268692   0.4244415760765611   0.9759013288431809   0.4458659959736642   0.26948923038135797   0.5710105035732242   0.08981732200385083   0.2941943510890242   0.8713619316138568   0.9108018458476497   0.5741389872314402   0.3428103024068045   0.02811383469506343   0.6904729092370258   0.8619948351091075   0.8700711806102215   0.3578967476940223   0.5371482717756382   0.3108536282761608   0.8191075383265402   0.3800240254504492   0.7178895636952547   0.7449157018650475   0.18221459077031588   0.2337007542877623   0.29344798761869356
0.7690143730218666   0.7363485947966516   0.9642115239064043   0.7224374840454694   0.6791970510180158   0.44215424370762746   0.09284959229254756   0.8116356381978196   0.10505806378657559   0.09934394130082295   0.06473575759748414   0.12116272896079383   0.24306322867746813   0.22927276069060146   0.7068390099034618   0.5840144571851557   0.9322096004013073   0.41016522236406133   0.3268149844530126   0.866124893489901   0.18729389853625977   0.22795063159374548   0.09311423016525026   0.5726769058712073   0.4182795255143932   0.49160203679709386   0.12890270625884592   0.8502394218257381   0.7390824744963774   0.04944779308946637   0.03605311396629836   0.03860378362791843   0.6340244107098019   0.9501038517886434   0.9713173563688142   0.9174410546671246   0.3909611820323337   0.720831091098042   0.2644783464653524   0.333426597481969   0.4587515816310264   0.3106658687339806   0.9376633620123398   0.46730170399206805   0.27145768309476664   0.08271523714023514   0.8445491318470896   0.8946247981208607   0.8531781575803734   0.5911132003431413   0.7156464255882437   0.04438537629512259   0.11409568308399605   0.541665407253675   0.6795933116219453   0.0057815926672041655   0.4800712723741942   0.5915615554650315   0.708275955253131   0.08834053800007957   0.08911009034186049   0.8707304643669895   0.44379760878777863   0.7549139405181106
0.6303585087108341   0.5600645956330089   0.5061342467754388   0.28761223652604256   0.35890082561606745   0.4773493584927738   0.6615851149283493   0.3929874384051819   0.505722668035694   0.8862361581496325   0.9459386893401056   0.3486020621100593   0.3916269849516979   0.34457075089595757   0.2663453777181603   0.34282046944285516   0.9115557125775037   0.753009195430926   0.5580694224650292   0.2544799314427756   0.8224456222356432   0.8822787310639365   0.11427181367725062   0.49956599092466497   0.19208711352480914   0.32221413543092753   0.6081375669018118   0.21195375439862243   0.8331862879087417   0.8448647769381538   0.9465524519734626   0.8189663159934405   0.32746361987304773   0.9586286187885212   0.0006137626333569562   0.47036425388338127   0.9358366349213498   0.6140578678925637   0.7342683849151966   0.1275437844405261   0.02428092234384611   0.8610486724616376   0.17619896245016736   0.8730638529977506   0.2018353001082029   0.9787699413977012   0.06192714877291675   0.37349786207308555   0.009748186583393735   0.6565558059667737   0.45378958187110496   0.16154410767446314   0.17656189867465202   0.8116910290286199   0.5072371298976424   0.3425777916810226   0.8490982788016043   0.8530624102400987   0.5066233672642855   0.8722135377976413   0.9132616438802544   0.23900454234753493   0.7723549823490888   0.7446697533571152
0.8889807215364083   0.37795586988589724   0.5961560198989214   0.8716059003593647   0.6871454214282054   0.39918592848819606   0.5342288711260047   0.4981080382862791   0.6773972348448117   0.7426301225214225   0.08043928925489972   0.33656393061181594   0.5008353361701597   0.9309390934928026   0.5732021593572574   0.9939861389307934   0.6517370573685555   0.07787668325270389   0.0665787920929719   0.12177260113315203   0.738475413488301   0.8388721409051689   0.2942238097438831   0.3771028477760368   0.8494946919518926   0.4609162710192717   0.6980677898449617   0.5054969474166722   0.1623492705236872   0.061730342531075615   0.16383891871895703   0.007388909130393082   0.4849520356788755   0.31910022000965316   0.0833996294640573   0.6708249785185771   0.9841166995087158   0.38816112651685064   0.5101974701067999   0.6768388395877838   0.33237964214016036   0.3102844432641467   0.44361867801382804   0.5550662384546318   0.5939042286518594   0.4714123023589778   0.14939486826994494   0.17796339067859493   0.7444095366999668   0.010496031339706098   0.45132707842498326   0.6724664432619227   0.5820602661762795   0.9487656888086304   0.2874881597060262   0.6650775341315297   0.09710823049740404   0.6296654687989773   0.20408853024196894   0.9942525556129526   0.11299153098868825   0.24150434228212667   0.693891060135169   0.31741371602516877
0.7806118888485278   0.93121989901798   0.2502723821213409   0.762347477570537   0.18670766019666848   0.4598075966590021   0.10087751385139598   0.5843840868919421   0.4422981234967017   0.44931156531929606   0.6495504354264128   0.9119176436300194   0.8602378573204222   0.5005458765106655   0.3620622757203865   0.24684010949848964   0.7631296268230182   0.8708804077116883   0.15797374547841755   0.2525875538855371   0.6501380958343299   0.6293760654295616   0.4640826853432486   0.9351738378603683   0.8695262069858021   0.6981561664115816   0.21381030322190767   0.17282636028983128   0.6828185467891336   0.2383485697525795   0.1129327893705117   0.5884422733978892   0.2405204232924318   0.7890370044332835   0.463382353944099   0.6765246297678699   0.3802825659720096   0.28849112792261794   0.10132007822371247   0.4296845202693802   0.6171529391489915   0.4176107202109297   0.9433463327452949   0.17709696638384312   0.9670148433146616   0.7882346547813681   0.4792636474020463   0.2419231285234748   0.09748863632885948   0.09007848836978648   0.26545334418013866   0.06909676823364352   0.41467008953972595   0.8517299186172069   0.15252055480962695   0.48065449483575434   0.1741496662472941   0.06269291418392346   0.689138200865528   0.8041298650678844   0.7938671002752845   0.7742017862613055   0.5878181226418155   0.3744453447985042
0.17671416112629304   0.3565910660503758   0.6444717898965205   0.1973483784146611   0.20969931781163148   0.5683564112690077   0.16520814249447427   0.9554252498911863   0.112210681482772   0.4782779228992212   0.8997547983143356   0.8863284816575427   0.6975405919430461   0.6265480042820143   0.7472342435047087   0.40567398682178846   0.523390925695752   0.5638550900980908   0.05809604263918071   0.601544121753904   0.7295238254204675   0.7896533038367852   0.47027791999736523   0.22709877695539976   0.5528096642941744   0.43306223778640945   0.8258061301008447   0.02975039854073865   0.34311034648254296   0.8647058265174018   0.6605979876063703   0.07432514864955236   0.23089966499977096   0.3864279036181805   0.7608431892920348   0.1879966669920096   0.5333590730567249   0.7598798993361663   0.013608945787326089   0.7823226801702211   0.00996814736097291   0.19602480923807547   0.9555129031481454   0.18077855841631715   0.28044432194050545   0.4063715054012902   0.4852349831507802   0.9536797814609174   0.727634657646331   0.9733092676148808   0.6594288530499355   0.9239293829201788   0.384524311163788   0.10860344109747899   0.9988308654435651   0.8496042342706264   0.15362464616401705   0.7221755374792984   0.23798767615153038   0.6616075672786168   0.6202655731072921   0.9622956381431322   0.2243787303642043   0.8792848871083957
0.6102974257463193   0.7662708289050567   0.2688658272160589   0.6985063286920785   0.32985310380581384   0.3598993235037666   0.7836308440652787   0.744826547231161   0.6022184461594828   0.38659005588888584   0.12420199101534322   0.8208971643109824   0.21769413499569484   0.27798661479140685   0.12537112557177807   0.9712929300403559   0.06406948883167779   0.5558110773121083   0.8873834494202477   0.3096853627617391   0.4438039157243856   0.5935154391689762   0.6630047190560434   0.43040047565334344   0.8335064899780663   0.8272446102639194   0.39413889183998446   0.731894146961265   0.5036533861722525   0.46734528676015286   0.6105080477747057   0.9870675997301038   0.9014349400127696   0.08075523087126701   0.4863060567593625   0.16617043541912152   0.6837408050170748   0.8027686160798602   0.36093493118758446   0.1948775053787656   0.619671316185397   0.2469575387677518   0.47355148176733675   0.8851921426170265   0.17586740046101138   0.6534420995987756   0.8105467627112933   0.45479166696368306   0.34236091048294504   0.8261974893348563   0.41640787087130887   0.7228975200024181   0.8387075243106925   0.3588522025747034   0.8058998230966031   0.7358299202723143   0.9372725842979229   0.2780969717034364   0.3195937663372406   0.5696594848531927   0.25353177928084814   0.4753283556235762   0.9586588351496561   0.37478197947442715
0.6338604630954511   0.22837081685582442   0.4851073533823194   0.48958983685740065   0.4579930626344398   0.5749287172570487   0.674560590671026   0.03479816989371758   0.11563215215149475   0.7487312279221925   0.2581527197997172   0.31190064989129945   0.27692462784080224   0.3898790253474891   0.4522528967031141   0.5760707296189852   0.33965204354287937   0.11178205364405269   0.13265913036587348   0.006411244765792374   0.08612026426203125   0.6364536980204765   0.17400029521621732   0.6316292652913652   0.4522598011665801   0.4080828811646521   0.6888929418338979   0.14203942843396455   0.9942667385321403   0.8331541639076033   0.014332351162871846   0.10724125854024696   0.8786345863806456   0.08442293598541079   0.7561796313631546   0.7953406086489475   0.6017099585398433   0.6945439106379216   0.30392673466004055   0.2192698790299624   0.262057914996964   0.582761856993869   0.17126760429416704   0.21285863426417   0.17593765073493275   0.9463081589733925   0.9972673090779497   0.5812293689728047   0.7236778495683527   0.5382252778087405   0.3083743672440518   0.43918994053884025   0.7294111110362123   0.7050711139011372   0.29404201608117997   0.3319486819985933   0.8507765246555667   0.6206481779157264   0.5378623847180253   0.5366080733496458   0.24906656611572334   0.9261042672778047   0.23393565005798478   0.31733819431968335
0.9870086511187594   0.34334241028393575   0.06266804576381772   0.10447956005551336   0.8110710003838265   0.3970342513105432   0.06540073668586802   0.5232501910827085   0.0873931508154739   0.8588089735018027   0.7570263694418162   0.08406025054386831   0.35798203977926163   0.15373785960066555   0.46298435336063626   0.752111568545275   0.5072055151236949   0.5330896816849392   0.925121968642611   0.2155034951956293   0.2581389490079716   0.6069854144071345   0.6911863185846262   0.8981653008759459   0.2711302978892123   0.26364300412319874   0.6285182728208084   0.7936857408204325   0.4600592975053857   0.8666087528126555   0.5631175361349404   0.270435549737724   0.3726661466899118   0.0077997793108527756   0.8060911666931242   0.1863752991938557   0.014684106910650203   0.8540619197101872   0.34310681333248794   0.43426373064858065   0.5074785917869553   0.32097223802524805   0.41798484468987696   0.21876023545295134   0.24933964277898368   0.7139868236181136   0.7267985261052508   0.32059493457700544   0.9782093448897714   0.45034381949491487   0.09828025328444231   0.5269091937565729   0.5181500473843857   0.5837350666822594   0.5351627171495019   0.2564736440188488   0.1454839006944739   0.5759352873714065   0.7290715504563776   0.07009834482499314   0.13079979378382367   0.7218733676612193   0.3859647371238897   0.6358346141764125
0.6233212019968684   0.4009011296359713   0.9679798924340127   0.41707437872346115   0.3739815592178847   0.6869143060178577   0.24118136632876194   0.09647944414645572   0.39577221432811327   0.23657048652294285   0.14290111304431963   0.5695702503898828   0.8776221669437276   0.6528354198406835   0.6077383958948178   0.31309660637103404   0.7321382662492537   0.07690013246927689   0.8786668454384401   0.2429982615460409   0.60133847246543   0.3550267648080575   0.4927021083145504   0.6071636473696284   0.9780172704685617   0.9541256351720862   0.5247222158805377   0.19008926864616726   0.6040357112506769   0.26721132915422846   0.2835408495517757   0.09360982449971154   0.20826349692256366   0.030640842631285626   0.1406397365074561   0.5240395741098287   0.33064132997883605   0.37780542279060214   0.5329013406126383   0.21094296773879465   0.5985030637295824   0.30090529032132524   0.6542344951741982   0.9679447061927537   0.9971645912641524   0.9458785255132677   0.16153238685964777   0.36078105882312533   0.0191473207955907   0.9917528903411815   0.6368101709791101   0.17069179017695807   0.4151116095449138   0.7245415611869531   0.35326932142733436   0.07708196567724653   0.20684811262235012   0.6939007185556675   0.21262958491987824   0.5530423915674179   0.876206782643514   0.3160952957650653   0.6797282443072399   0.3420994238286232
0.2777037189139317   0.015190005443740048   0.025493749133041716   0.37415471763586944   0.28053912764977934   0.06931147993047232   0.8639613622733939   0.013373658812744122   0.26139180685418867   0.07755858958929078   0.22715119129428385   0.8426818686357861   0.8462801973092748   0.35301702840233773   0.8738818698669495   0.7655999029585395   0.6394320846869248   0.6591163098466702   0.6612522849470712   0.2125575113911217   0.7632253020434108   0.34302101408160496   0.9815240406398313   0.8704580875624985   0.485521583129479   0.3278310086378649   0.9560302915067896   0.49630336992662905   0.20498245547969968   0.2585195287073926   0.0920689292333957   0.4829297111138849   0.943590648625511   0.18096093911810182   0.8649177379391119   0.6402478424780988   0.09731045131623613   0.8279439107157641   0.9910358680721624   0.8746479395195593   0.45787836662931136   0.16882760086909385   0.32978358312509104   0.6620904281284377   0.6946530645859006   0.8258065867874889   0.3482595424852597   0.7916323405659391   0.20913148145642158   0.49797557814962395   0.39222925097847006   0.29532897063931013   0.0041490259767218984   0.2394560494422313   0.30016032174507434   0.8123992595254252   0.060558377351210876   0.05849511032412949   0.4352425838059625   0.17215141704732634   0.9632479260349748   0.23055119960836537   0.44420671573380016   0.297503477527767
0.5053695594056634   0.061723598739271544   0.11442313260870912   0.6354130493993294   0.8107164948197627   0.2359170119517827   0.7661635901234495   0.8437807088333903   0.6015850133633411   0.7379414338021587   0.3739343391449794   0.5484517381940801   0.5974359873866193   0.49848538435992745   0.07377401739990505   0.736052478668655   0.5368776100354085   0.43999027403579793   0.6385314335939426   0.5639010616213286   0.5736296840004337   0.20943907442743256   0.19432471786014238   0.26639758409356157   0.06826012459477028   0.147715475688161   0.07990158525143326   0.6309845346942322   0.2575436297750075   0.9117984637363783   0.31373799512798384   0.787203825860842   0.6559586164116663   0.1738570299342196   0.9398036559830044   0.23875208766676184   0.05852262902504705   0.6753716455742922   0.8660296385830993   0.502699608998107   0.5216450189896387   0.2353813715384942   0.22749820498915682   0.9387985473767783   0.948015334989205   0.02594229711106164   0.03317348712901443   0.6724009632832167   0.8797552103944347   0.8782268214229006   0.9532719018775812   0.04141642858898449   0.6222115806194272   0.9664283576865222   0.6395339067495973   0.2542126027281425   0.9662529642077609   0.7925713277523027   0.6997302507665929   0.015460515061380669   0.9077303351827138   0.11719968217801055   0.8337006121834936   0.5127609060632737
0.3860853161930751   0.8818183106395163   0.6062024071943367   0.5739623586864955   0.4380699812038702   0.8558760135284547   0.5730289200653222   0.9015613954032787   0.5583147708094355   0.9776491921055541   0.6197570181877411   0.8601449668142943   0.9361031901900083   0.011220834419031805   0.9802231114381438   0.6059323640861517   0.9698502259822475   0.2186495066667291   0.2804928606715509   0.5904718490247711   0.06211989079953369   0.10144982448871856   0.4467922484880573   0.07771094296149732   0.6760345746064585   0.2196315138492022   0.8405898412937206   0.5037485842750019   0.23796459340258835   0.3637555003207475   0.26756092122839825   0.6021871888717231   0.6796498225931529   0.38610630821519343   0.6478039030406572   0.7420422220574289   0.7435466324031446   0.3748854737961616   0.6675807916025134   0.1361098579712771   0.7736964064208971   0.15623596712943252   0.3870879309309625   0.545638008946506   0.7115765156213634   0.05478614264071395   0.9402956824429052   0.46792706598500866   0.03554194101490483   0.8351546287915117   0.09970584114918464   0.9641784817100069   0.7975773476123165   0.4713991284707642   0.8321449199207863   0.36199129283828374   0.1179275250191636   0.08529282025557079   0.18434101688012922   0.6199490707808549   0.37438089261601903   0.7104073464594092   0.5167602252776159   0.4838392128095778
0.6006844861951219   0.5541713793299766   0.12967229434665334   0.9382012038630718   0.8891079705737586   0.4993852366892627   0.1893766119037481   0.4702741378780631   0.8535660295588537   0.664230607897751   0.08967077075456348   0.5060956561680563   0.05598868194653732   0.19283147942698675   0.2575258508337771   0.14410436332977256   0.9380611569273737   0.10753865917141595   0.07318483395364789   0.5241552925489177   0.5636802643113547   0.3971313127120068   0.556424608676032   0.04031607973933985   0.9629957781162327   0.8429599333820301   0.4267523143293787   0.10211487587626804   0.07388780754247407   0.3435746966927674   0.2373757024256306   0.631840737998205   0.22032177798362026   0.6793440887950164   0.14770493167106713   0.12574508183014863   0.16433309603708296   0.4865126093680297   0.89017908083729   0.981640718500376   0.22627193910970922   0.37897395019661373   0.8169942468836421   0.4574854259514584   0.6625916747983546   0.981842637484607   0.2605696382076101   0.41716934621211854   0.6995958966821219   0.13888270410257686   0.8338173238782314   0.3150544703358505   0.6257080891396478   0.7953080074098094   0.5964416214526007   0.6832137323376456   0.4053863111560276   0.11596391861479301   0.44873668978153364   0.5574686505074969   0.24105321511894462   0.6294513092467633   0.5585576089442437   0.5758279320071209
0.014781276009235372   0.25047735905014956   0.7415633620606015   0.11834250605566249   0.35218960121088083   0.26863472156554263   0.48099372385299144   0.7011731598435439   0.6525937045287589   0.12975201746296577   0.6471763999747601   0.38611868950769346   0.02688561538911109   0.3344440100531563   0.05073477852215934   0.7029049571700479   0.6214993042330835   0.2184800914383633   0.6019980887406257   0.14543630666255092   0.3804460891141389   0.5890287821915999   0.04344047979638208   0.56960837465543   0.36566481310490356   0.33855142314145037   0.3018771177357806   0.45126586859976753   0.013475211894022744   0.06991670157590778   0.8208833938827891   0.7500927087562236   0.3608815073652638   0.940164684112942   0.17370699390802904   0.3639740192485301   0.33399589197615276   0.6057206740597857   0.12297221538586971   0.6610690620784823   0.7124965877430692   0.3872405826214224   0.520974126645244   0.5156327554159313   0.33205049862893027   0.7982118004298224   0.4775336468488619   0.9460243807605013   0.9663856855240267   0.45966037728837206   0.17565652911308133   0.4947585121607338   0.952910473630004   0.38974367571246427   0.3547731352302922   0.7446658034045103   0.5920289662647402   0.44957899159952225   0.18106614132226315   0.3806917841559801   0.2580330742885874   0.8438583175397365   0.058093925936393453   0.7196227220774978
0.5455364865455182   0.45661773491831414   0.5371197992911495   0.2039899666615664   0.21348598791658793   0.6584059344884917   0.05958615244228756   0.25796558590106505   0.2471003023925612   0.1987455572001197   0.8839296233292062   0.7632070737403313   0.2941898287625572   0.8090018814876554   0.529156488098914   0.018541270335821005   0.7021608624978171   0.3594228898881332   0.34809034677665085   0.6378494861798409   0.4441277882092296   0.5155645723483966   0.2899964208402574   0.9182267641023432   0.8985913016637114   0.05894683743008249   0.752876621549108   0.7142367974407767   0.6851053137471235   0.4005409029415908   0.6932904691068204   0.4562712115397117   0.43800501135456227   0.20179534574147107   0.8093608457776141   0.6930641377993805   0.14381518259200507   0.3927934642538156   0.28020435767870017   0.6745228674635594   0.44165432009418804   0.03337057436568245   0.9321140109020493   0.0366733812837185   0.9975265318849584   0.5178060020172858   0.6421175900617918   0.11844661718137536   0.09893523022124703   0.4588591645872033   0.8892409685126839   0.40420981974059866   0.4138299164741236   0.05831826164561255   0.19595049940586348   0.9479386082008869   0.9758249051195613   0.8565229159041415   0.3865896536282493   0.2548744704015065   0.8320097225275562   0.46372945165032586   0.10638529594954917   0.5803516029379471
0.3903554024333682   0.4303588772846434   0.1742712850474999   0.5436782216542286   0.39282887054840976   0.9125528752673576   0.5321536949857081   0.42523160447285324   0.2938936403271627   0.4536937106801543   0.6429127264730242   0.02102178473225461   0.8800637238530391   0.3953754490345417   0.4469622270671607   0.07308317653136763   0.9042388187334779   0.5388525331304003   0.06037257343891138   0.8182087061298611   0.07222909620592162   0.07512308148007439   0.9539872774893622   0.23785710319191397   0.6818736937725535   0.644764204195431   0.7797159924418623   0.6941788815376854   0.2890448232241437   0.7322113289280734   0.24756229745615424   0.2689472770648321   0.995151182896981   0.27851761824791915   0.6046495709831301   0.24792549233257752   0.11508745904394187   0.8831421692133774   0.1576873439159694   0.17484231580120987   0.21084864031046402   0.3442896360829772   0.097314770477058   0.3566336096713488   0.13861954410454239   0.2691665546029028   0.1433274929876958   0.1187765064794348   0.45674585033198895   0.6244023504074718   0.36361150054583347   0.42459762494174946   0.16770102710784524   0.8921910214793984   0.11604920308967923   0.1556503478769173   0.17254984421086425   0.6136734032314792   0.5113996321065492   0.9077248555443398   0.057462385166922376   0.7305312340181018   0.35371228819057976   0.7328825397431299
0.8466137448564584   0.38624159793512464   0.25639751771352176   0.3762489300717812   0.707994200751916   0.11707504333222184   0.11307002472582597   0.25747242359234634   0.251248350419927   0.49267269292475   0.7494585241799925   0.8328747986505969   0.08354732331208176   0.6004816714453516   0.6334093210903132   0.6772244507736797   0.9109974791012175   0.9868082682138724   0.12200968898376412   0.7694995952293398   0.8535350939342952   0.2562770341957705   0.7682974007931843   0.036617055486209846   0.006921349077836789   0.8700354362606458   0.5118998830796626   0.6603681254144287   0.2989271483259208   0.752960392928424   0.3988298583538366   0.40289570182208234   0.04767879790599383   0.260287700003674   0.6493713341738441   0.5700209031714853   0.964131474593912   0.6598060285583224   0.01596201308353084   0.8927964523978058   0.05313399549269455   0.67299776034445   0.8939523240997668   0.12329685716846601   0.1995989015583994   0.4167207261486795   0.12565492330658237   0.08667980168225617   0.19267755248056262   0.5466852898880337   0.6137550402269198   0.42631167626782746   0.8937504041546418   0.7937248969596096   0.2149251818730832   0.02341597444574515   0.846071606248648   0.5334371969559356   0.5655538476992391   0.45339507127425976   0.8819401316547358   0.8736311683976132   0.5495918346157083   0.5605986188764539
0.8288061361620414   0.20063340805316315   0.6556395105159415   0.43730176170798796   0.6292072346036419   0.7839126819044837   0.5299845872093591   0.35062196002573176   0.4365296821230793   0.23722739201645004   0.9162295469824393   0.9243102837579042   0.5427792779684375   0.4435024950568404   0.7013043651093561   0.9008943093121592   0.6967076717197895   0.9100652981009049   0.13575051741011704   0.44749923803789937   0.8147675400650537   0.036434129703291664   0.5861586827944087   0.8869006191614455   0.9859614039030123   0.8358007216501285   0.9305191722784673   0.4495988574534575   0.3567541692993704   0.051888039745644834   0.40053458506910805   0.09897689742772574   0.9202244871762911   0.8146606477291948   0.48430503808666875   0.17466661366982145   0.3774452092078536   0.37115815267235436   0.7830006729773126   0.2737723043576623   0.680737537488064   0.4610928545714495   0.6472501555671956   0.8262730663197629   0.8659699974230104   0.4246587248681578   0.0610914727727868   0.9393724471583175   0.880008593519998   0.5888580032180293   0.1305723004943196   0.48977358970485996   0.5232544242206275   0.5369699634723845   0.7300377154252115   0.3907966922771342   0.6030299370443365   0.7223093157431897   0.24573267733854276   0.21613007860731276   0.22558472783648284   0.3511511630708353   0.4627320043612302   0.9423577742496504
0.5448471903484188   0.8900583084993858   0.8154818487940346   0.11608470792988752   0.6788771929254085   0.465399583631228   0.7543903760212478   0.17671226077157007   0.7988685994054104   0.8765415804131986   0.6238180755269283   0.6869386710667101   0.2756141751847829   0.33957161694081417   0.8937803601017167   0.2961419787895759   0.6725842381404464   0.6172623011976245   0.6480476827631739   0.08001190018226313   0.4469995103039636   0.26611113812678916   0.1853156784019438   0.1376541259326127   0.9021523199555448   0.37605282962740333   0.36983382960790917   0.021569418002725157   0.22327512703013636   0.9106532459961753   0.6154434535866614   0.8448571572311551   0.4244065276247259   0.034111665582976645   0.9916253780597332   0.15791848616444498   0.14879235243994302   0.6945400486421625   0.09784501795801641   0.8617765073748691   0.47620811429949655   0.07727774744453801   0.44979733519484244   0.781764607192606   0.029208603995532958   0.8111666093177489   0.26448165679289865   0.6441104812599933   0.12705628403998814   0.4351137796903456   0.8946478271849895   0.6225410632572681   0.9037811570098518   0.5244605336941702   0.2792043735983281   0.777683906026113   0.47937462938512587   0.4903488681111936   0.28757899553859495   0.619765419861668   0.3305822769451829   0.7958088194690311   0.18973397758057856   0.7579889124867989
0.8543741626456863   0.7185310720244932   0.7399366423857361   0.976224305294193   0.8251655586501534   0.9073644627067442   0.47545498559283744   0.3321138240341997   0.6981092746101653   0.47225068301639866   0.580807158407848   0.7095727607769315   0.7943281176003134   0.9477901493222284   0.3016027848095199   0.9318888547508185   0.31495348821518754   0.4574412812110348   0.01402378927092493   0.31212343488915045   0.9843712112700046   0.6616324617420036   0.8242898116903464   0.5541345224023515   0.12999704862431832   0.9431013897175106   0.08435316930461027   0.5779102171081586   0.304831489974165   0.035736927010766265   0.6088981837117728   0.2457963930739589   0.6067222153639997   0.5634862439943676   0.02809102530392483   0.5362236322970273   0.8123940977636863   0.6156960946721391   0.726488240494405   0.6043347775462088   0.49744060954849884   0.15825481346110443   0.71246445122348   0.29221134265705834   0.5130693982784942   0.4966223517191008   0.8881746395331336   0.7380768202547068   0.3830723496541759   0.5535209620015903   0.8038214702285233   0.16016660314654824   0.07824085968001092   0.517784034990824   0.19492328651675053   0.9143702100725893   0.47151864431601115   0.9542977909964564   0.1668322612128257   0.378146577775562   0.6591245465523248   0.3386016963243172   0.44034402071842077   0.7738118002293531
0.16168393700382594   0.1803468828632128   0.7278795694949408   0.4816004575722948   0.6486145387253317   0.683724531144112   0.8397049299618071   0.743523637317588   0.26554218907115584   0.1302035691425217   0.035883459733283773   0.5833570341710398   0.18730132939114494   0.6124195341516977   0.8409601732165333   0.6689868240984504   0.7157826850751338   0.6581217431552413   0.6741279120037075   0.2908402463228884   0.05665813852280898   0.31952004683092405   0.23378389128528673   0.5170284460935353   0.894974201518983   0.1391731639677113   0.505904321790346   0.035427988521240406   0.2463596627936513   0.4554486328235993   0.6661993918285388   0.2919043512036524   0.9808174737224954   0.3252450636810776   0.630315932095255   0.7085473170326126   0.7935161443313505   0.7128255295293798   0.7893557588787218   0.0395604929341622   0.07773345925621675   0.05470378637413859   0.11522784687501432   0.7487202466112738   0.021075320733407763   0.7351837395432145   0.8814439555897275   0.23169180051773855   0.12610111921442474   0.5960105755755032   0.3755396337993816   0.19626381199649814   0.8797414564207734   0.14056194275190392   0.7093402419708428   0.9043594607928458   0.898923982698278   0.8153168790708263   0.0790243098755877   0.19581214376023312   0.10540783836692748   0.10249134954144645   0.2896685509968659   0.15625165082607093
0.02767437911071073   0.04778756316730785   0.17444070412185156   0.4075314042147971   0.006599058377302966   0.31260382362409334   0.292996748532124   0.1758396036970586   0.8804979391628782   0.7165932480485901   0.9174571147327424   0.9795757917005604   0.000756482742104796   0.5760313052966862   0.20811687276189964   0.07521633090771467   0.10183250004382681   0.7607144262258598   0.12909256288631193   0.8794041871474816   0.9964246616768994   0.6582230766844134   0.839424011889446   0.7231525363214106   0.9687502825661886   0.6104355135171056   0.6649833077675945   0.31562113210661347   0.9621512241888857   0.29783168989301223   0.3719865592354705   0.1397815284095549   0.0816532850260074   0.5812384418444221   0.45452944450272814   0.16020573670899446   0.0808968022839026   0.005207136547735908   0.2464125717408285   0.0849894058012798   0.9790643022400758   0.24449271032187606   0.11732000885451657   0.20558521865379825   0.9826396405631764   0.5862696336374627   0.2778959969650705   0.4824326823323877   0.013889357996987869   0.9758341201203571   0.612912689197476   0.16681155022577418   0.05173813380810224   0.6780024302273449   0.24092612996200552   0.027030021816219277   0.9700848487820949   0.09676398838292273   0.7863966854592774   0.8668242851072248   0.8891880464981923   0.09155685183518683   0.5399841137184489   0.781834879305945
0.9101237442581165   0.8470641415133108   0.4226641048639323   0.5762496606521468   0.9274841036949399   0.2607945078758482   0.1447681078988618   0.09381697831975909   0.9135947456979521   0.2849603877554911   0.5318554187013858   0.9270054280939849   0.8618566118898499   0.6069579575281463   0.29092928873938023   0.8999754062777656   0.8917717631077551   0.5101939691452235   0.5045326032801029   0.03315112117054083   0.002583716609562788   0.41863711731003667   0.964548489561654   0.25131624186459584   0.09245997235144635   0.571572975796726   0.5418843846977217   0.6750665812124491   0.16497586865650637   0.31077846792087777   0.3971162767988599   0.58124960289269   0.25138112295855425   0.02581808016538666   0.8652608580974741   0.6542441747987051   0.3895245110687044   0.41886012263724043   0.5743315693580939   0.7542687685209395   0.49775274796094937   0.9086661534920168   0.06979896607799102   0.7211176473503986   0.49516903135138657   0.4900290361819802   0.10525047651633702   0.4698014054858028   0.40270905899994025   0.9184560603852543   0.5633660918186153   0.7947348242733537   0.23773319034343388   0.6076775924643766   0.16624981501975544   0.21348522138066373   0.9863520673848796   0.5818595122989899   0.30098895692228134   0.5592410465819586   0.5968275563161752   0.16299938966174948   0.7266573875641874   0.8049722780610192
0.09907480835522581   0.2543332361697326   0.6568584214861964   0.08385463071062059   0.6039057770038392   0.7643041999877523   0.5516079449698594   0.6140532252248178   0.201196718003899   0.845848139602498   0.988241853151244   0.8193184009514641   0.9634635276604651   0.23817054713812152   0.8219920381314886   0.6058331795708004   0.9771114602755855   0.6563110348391317   0.5210030812092072   0.04659213298884172   0.3802839039594103   0.4933116451773822   0.7943456936450198   0.2416198549278225   0.2812090956041845   0.2389784090076496   0.13748727215882345   0.15776522421720193   0.6773033186003453   0.4746742090198972   0.5858793271889641   0.5437119989923841   0.4761066005964463   0.6288260694173992   0.59763747403772   0.7243935980409201   0.5126430729359812   0.39065552227927763   0.7756454359062315   0.11856041847011968   0.5355316126603957   0.7343444874401459   0.2546423546970241   0.07196828548127795   0.15524770870098537   0.24103284226276378   0.4602966610520043   0.8303484305534554   0.8740386130968009   0.00205443325511419   0.32280938889318084   0.6725832063362536   0.19673529449645558   0.527380224235217   0.7369300617042167   0.1288712073438694   0.7206286939000093   0.8985541548178179   0.13929258766649674   0.40447760930294935   0.20798562096402806   0.5078986325385402   0.3636471517602653   0.2859171908328297
0.6724540083036323   0.7735541450983943   0.10900479706324119   0.21394890535155173   0.517206299602647   0.5325213028356305   0.6487081360112369   0.3836004747980963   0.6431676865058461   0.5304668695805163   0.3258987471180561   0.7110172684618428   0.44643239200939056   0.003086645345299303   0.5889686854138394   0.5821460611179734   0.7258036981093813   0.10453249052748148   0.44967609774734263   0.177668451815024   0.5178180771453532   0.5966338579889413   0.0860289459870773   0.8917512609821943   0.8453640688417209   0.823079712890547   0.9770241489238362   0.6778023556306426   0.32815776923907386   0.29055841005491656   0.3283160129125992   0.29420188083254634   0.6849900827332277   0.7600915404744003   0.00241726579454308   0.5831846123707036   0.23855769072383715   0.757004895129101   0.4134485803807037   0.0010385512527302345   0.5127539926144559   0.6524724046016195   0.9637724826333611   0.8233700994377062   0.9949359154691026   0.05583854661267824   0.8777435366462838   0.931618838455512   0.14957184662738177   0.23275883372213121   0.9007193877224476   0.25381648282486935   0.821414077388308   0.9422004236672147   0.5724033748098485   0.9596146019923231   0.13642399465508023   0.18210888319281437   0.5699861090153054   0.37642998962161944   0.8978663039312431   0.42510398806371336   0.15653752863460169   0.3753914383688892
0.38511231131678725   0.7726315834620938   0.1927650460012406   0.552021338931183   0.39017639584768465   0.7167930368494156   0.31502150935495676   0.620402500475671   0.24060454922030286   0.4840342031272844   0.4143021216325091   0.3665860176508017   0.4191904718319949   0.5418337794600697   0.8418987468226606   0.40697141565847866   0.28276647717691467   0.3597248962672554   0.2719126378073552   0.030541426036859227   0.3849001732456716   0.934620908203542   0.11537510917275348   0.6551499876679701   0.9997878619288844   0.16198932474144817   0.9226100631715128   0.10312864873678707   0.6096114660811996   0.4451962878920325   0.6075885538165561   0.48272614826111604   0.3690069168608968   0.9611620847647482   0.193286432184047   0.11614013061031438   0.949816445028902   0.41932830530467835   0.3513876853613864   0.7091687149518358   0.6670499678519872   0.05960340903742298   0.07947504755403122   0.6786272889149765   0.2821497946063157   0.12498250083388095   0.9640999383812777   0.023477301247006453   0.2823619326774313   0.9629931760924328   0.04148987520976485   0.9203486525102194   0.6727504665962316   0.5177968882004003   0.43390132139320875   0.4376225042491033   0.3037435497353348   0.5566348034356521   0.24061488920916174   0.32148237363878895   0.3539271047064329   0.13730649813097376   0.8892272038477753   0.6123136586869532
0.6868771368544456   0.07770308909355078   0.8097521562937441   0.9336863697719767   0.40472734224813   0.9527205882596699   0.8456522179124664   0.9102090685249703   0.12236540957069868   0.989727412167237   0.8041623427027015   0.9898604160147509   0.449614942974467   0.47193052396683677   0.3702610213094928   0.5522379117656476   0.14587139323913226   0.9152957205311847   0.12964613210033105   0.23075553812685864   0.7919442885326994   0.7779892224002108   0.2404189282525557   0.6184418794399054   0.10506715167825371   0.7002861333066601   0.4306667719588116   0.6847555096679286   0.7003398094301237   0.7475655450469902   0.5850145540463452   0.7745464411429583   0.577974399859425   0.7578381328797532   0.7808522113436437   0.7846860251282074   0.128359456884958   0.28590760891291644   0.4105911900341509   0.23244811336255977   0.9824880636458257   0.3706118883817318   0.28094505793381985   0.001692575235701126   0.19054377511312637   0.5926226659815209   0.04052612968126412   0.38325069579579574   0.08547662343487265   0.8923365326748608   0.6098593577224526   0.6984951861278671   0.3851368140047489   0.14477098762787052   0.02484480367610734   0.9239487449849088   0.8071624141453239   0.3869328547481173   0.24399259233246368   0.13926271985670138   0.6788029572603659   0.10102524583520082   0.8334014022983128   0.9068146064941416
0.6963148936145401   0.730413357453469   0.552456344364493   0.9051220312584405   0.5057711185014138   0.1377906914719481   0.5119302146832289   0.5218713354626447   0.42029449506654115   0.24545415879708732   0.9020708569607763   0.8233761493347777   0.0351576810617922   0.1006831711692168   0.877226053284669   0.8994274043498689   0.2279952669164683   0.7137503164210995   0.6332334609522053   0.7601646844931675   0.5491923096561024   0.6127250705858988   0.7998320586538925   0.853350077999026   0.8528774160415623   0.8823117131324297   0.24737571428939953   0.9482280467405855   0.3471062975401485   0.7445210216604816   0.7354454996061707   0.42635671127794067   0.9268118024736074   0.49906686286339424   0.8333746426453944   0.602980561943163   0.8916541214118151   0.3983836916941775   0.9561485893607254   0.7035531575932941   0.6636588544953468   0.684633375273078   0.32291512840852016   0.9433884731001266   0.11446654483924443   0.07190830468717925   0.5230830697546276   0.09003839510110068   0.2615891287976822   0.18959659155474956   0.2757073554652281   0.14181034836051523   0.9144828312575337   0.445075569894268   0.5402618558590574   0.7154536370825746   0.9876710287839263   0.9460087070308737   0.7068872132136631   0.11247307513941154   0.09601690737211122   0.5476250153366963   0.7507386238529377   0.40891991754611745
0.4323580528767644   0.8629916400636183   0.4278234954444175   0.4655314444459908   0.3178915080375199   0.791083335376439   0.9047404256897899   0.3754930493448902   0.056302379239837774   0.6014867438216895   0.6290330702245618   0.23368270098437494   0.14181954798230406   0.15641117392742152   0.0887712143655043   0.5182290639018003   0.15414851919837771   0.2104024668965478   0.38188400115184123   0.40575598876238883   0.05813161182626649   0.6627774515598516   0.6311453772989036   0.9968360712162714   0.6257735589495022   0.7997858114962333   0.20332188185448613   0.5313046267702806   0.3078820509119822   0.008702476119794227   0.2985814561646963   0.1558115774253904   0.2515796716721444   0.40721573229810476   0.6695483859401345   0.9221288764410155   0.10976012368984032   0.2508045583706832   0.5807771715746303   0.4038998125392151   0.9556116044914627   0.040402091474135426   0.198893170422789   0.9981438237768262   0.8974799926651962   0.37762463991428386   0.5677477931238853   0.0013077525605548214   0.27170643371569403   0.5778388284180506   0.36442591126939927   0.47000312579027426   0.9638243828037119   0.5691363522982563   0.06584445510470298   0.31419154836488383   0.7122447111315674   0.16192062000015162   0.39629606916456844   0.3920626719238684   0.6024845874417272   0.9111160616294683   0.8155188975899382   0.9881628593846533
0.6468729829502645   0.8707139701553329   0.6166257271671491   0.9900190356078271   0.7493929902850683   0.4930893302410491   0.0488779340432638   0.9887112830472723   0.47768655656937437   0.9152505018229985   0.6844520227738645   0.518708157256998   0.5138621737656626   0.3461141495247422   0.6186075676691616   0.20451660889211415   0.8016174626340951   0.18419352952459053   0.2223114985045931   0.8124539369682457   0.19913287519236794   0.27307746789512216   0.40679260091465497   0.8242910775835924   0.5522598922421035   0.4023634977397892   0.7901668737475057   0.8342720419757654   0.802866901957035   0.90927416749874   0.7412889397042419   0.8455607589284931   0.32518034538766066   0.9940236656757415   0.05683691693037742   0.32685260167149516   0.8113181716219982   0.6479095161509993   0.4382293492612159   0.122335992779381   0.009700708987903093   0.46371598662640884   0.21591785075662273   0.3098820558111352   0.8105678337955351   0.19063851873128673   0.8091252498419678   0.48559097822754277   0.25830794155343173   0.7882750209914975   0.01895837609446204   0.6513189362517774   0.45544103959639665   0.8790008534927575   0.27766943639022007   0.8057581773232843   0.13026069420873598   0.884977187817016   0.22083251945984267   0.4789055756517891   0.31894252258673783   0.23706767166601653   0.7826031701986268   0.35656958287240814
0.30924181359883474   0.7733516850396076   0.5666853194420041   0.04668752706127289   0.4986739798032996   0.5827131663083209   0.7575600696000363   0.5610965488337302   0.24036603824986785   0.7944381453168234   0.7386016935055743   0.9097776125819528   0.7849249986534712   0.915437291824066   0.4609322571153541   0.1040194352586685   0.6546643044447352   0.030460104007050005   0.24009973765551149   0.6251138596068794   0.3357217818579974   0.7933924323410335   0.45749656745688466   0.2685442767344713   0.026479968259162667   0.02004074730142583   0.8908112480148807   0.22185674967319838   0.5278059884558631   0.43732758099310487   0.13325117841484435   0.6607602008394683   0.2874399502059952   0.6428894356762815   0.39464948490927015   0.7509825882575155   0.502514951552524   0.7274521438522156   0.933717227793916   0.646963152998847   0.8478506471077888   0.6969920398451656   0.6936174901384046   0.02184929339196763   0.5121288652497914   0.903599607504132   0.23612092268151985   0.7533050166574964   0.48564889699062874   0.8835588602027062   0.3453096746666392   0.5314482669842979   0.9578429085347657   0.4462312792096014   0.21205849625179488   0.8706880661448297   0.6704029583287704   0.8033418435333198   0.8174090113425247   0.11970547788731419   0.1678880067762464   0.07588969968110429   0.8836917835486087   0.4727423248884672
0.3200373596684576   0.3788976598359387   0.19007429341020418   0.45089303149649956   0.8079084944186662   0.4752980523318066   0.9539533707286844   0.6975880148390032   0.3222595974280374   0.5917391921291004   0.6086436960620452   0.16613974785470523   0.3644166888932717   0.14550791291949902   0.39658519981025026   0.2954516817098755   0.6940137305645012   0.34216606938617916   0.5791761884677256   0.17574620382256131   0.5261257237882548   0.26627636970507484   0.6954844049191168   0.7030038789340941   0.20608836411979728   0.8873787098691361   0.5054101115089127   0.2521108474375946   0.3981798697011311   0.41208065753732953   0.5514567407802283   0.5545228325985915   0.07592027227309375   0.8203414654082292   0.9428130447181832   0.3883830847438862   0.711503583379822   0.6748335524887301   0.546227844907933   0.0929314030340107   0.017489852815320804   0.332667483102551   0.9670516564402074   0.9171851992114494   0.49136412902706594   0.06639111339747611   0.2715672515210906   0.21418132027735523   0.2852757649072687   0.17901240352833994   0.7661571400121779   0.9620704728397607   0.8870958952061375   0.7669317459910104   0.2147003992319497   0.4075476402411692   0.8111756229330438   0.9465902805827813   0.2718873545137665   0.019164555497282975   0.09967203955322175   0.2717567280940511   0.7256595096058336   0.9262331524632723
0.08218218673790095   0.9390892449915001   0.7586078531656261   0.00904795325182287   0.590818057710835   0.872698131594024   0.4870406016445355   0.7948666329744676   0.3055422928035663   0.6936857280656841   0.7208834616323575   0.832796160134707   0.41844639759742874   0.9267539820746736   0.5061830624004078   0.4252485198935378   0.607270774664385   0.9801637014918924   0.2342957078866413   0.4060839643962548   0.5075987351111632   0.7084069733978413   0.5086361982808077   0.47985081193298257   0.4254165483732622   0.7693177284063412   0.7500283451151817   0.4708028586811597   0.8345984906624272   0.8966195968123171   0.2629877434706462   0.6759362257066921   0.5290561978588609   0.202933868746633   0.5421042818382887   0.8431400655719851   0.11060980026143219   0.27617988667195936   0.035921219437880895   0.4178915456784473   0.5033390255970472   0.29601618518006695   0.8016255115512396   0.011807581282192413   0.9957402904858841   0.5876092117822257   0.2929893132704318   0.5319567693492099   0.5703237421126218   0.8182914833758846   0.5429609681552502   0.061153910668050135   0.7357252514501946   0.9216718865635675   0.279973224684604   0.38521768496135805   0.20666905359133372   0.7187380178169345   0.7378689428463153   0.542077619389373   0.09605925332990153   0.44255813114497516   0.7019477234084344   0.12418607371092576
0.5927202277328543   0.1465419459649082   0.9003222118571949   0.11237849242873334   0.5969799372469702   0.5589327341826825   0.607332898586763   0.5804217230795234   0.026656195134348318   0.7406412508067979   0.06437193043151279   0.5192678124114734   0.2909309436841537   0.8189693642432304   0.7843987057469087   0.1340501274501153   0.08426189009281995   0.10023134642629586   0.04652976290059347   0.5919725080607423   0.9882026367629184   0.6576732152813207   0.34458203949215904   0.46778643434981654   0.39548240903006415   0.5111312693164125   0.44425982763496424   0.3554079419210832   0.798502471783094   0.95219853513373   0.8369269290482013   0.7749862188415597   0.7718462766487456   0.21155728432693216   0.7725549986166885   0.25571840643008636   0.48091533296459194   0.3925879200837018   0.9881562928697797   0.12166827897997105   0.396653442871772   0.2923565736574059   0.9416265299691862   0.5296957709192288   0.4084508061088536   0.6346833583760852   0.5970444904770271   0.06190933656941222   0.012968397078789473   0.1235520890596727   0.15278466284206293   0.7065013946483291   0.21446592529569553   0.17135355392594268   0.3158577337938617   0.9315151758067693   0.4426196486469499   0.9597962695990105   0.5433027351771732   0.675796769376683   0.9617043156823579   0.5672083495153087   0.5551464423073935   0.5541284903967119
0.565050872810586   0.2748517758579028   0.6135199123382072   0.024432719477483145   0.15660006670173235   0.6401684174818176   0.016475421861180117   0.9625233829080709   0.14363166962294288   0.5166163284221449   0.8636907590191172   0.25602198825974193   0.9291657443272473   0.34526277449620224   0.5478330252252556   0.3245068124529726   0.48654609568029744   0.3854665048971917   0.004530290048082348   0.6487100430762897   0.5248417799979395   0.818258155381883   0.44938384774068885   0.09458155267957773   0.9597909071873535   0.5434063795239802   0.8358639354024816   0.07014883320209458   0.8031908404856212   0.9032379620421626   0.8193885135413015   0.10762545029402366   0.6595591708626783   0.38662163362001767   0.9556977545221843   0.8516034620342817   0.7303934265354309   0.041358859123815414   0.40786472929692874   0.5270966495813092   0.24384733085513352   0.6558923542266237   0.4033344392488464   0.8783866065050195   0.7190055508571941   0.8376341988447408   0.9539505915081575   0.7838050538254417   0.7592146436698405   0.2942278193207606   0.11808665610567595   0.7136562206233472   0.9560238031842193   0.39098985727859803   0.2986981425643745   0.6060307703293235   0.296464632321541   0.00436822365858037   0.34300038804219024   0.7544273082950418   0.5660712057861101   0.9630093645347649   0.9351356587452615   0.22733065871373265
0.3222238749309766   0.30711701030814126   0.5318012194964151   0.3489440522087131   0.6032183240737825   0.46948281146340054   0.5778506279882576   0.5651389983832713   0.844003680403942   0.17525499214263998   0.45976397188258167   0.8514827777599242   0.8879798772197227   0.7842651348640419   0.16106582931820718   0.24545200743060064   0.5915152448981816   0.7798969112054616   0.818065441276017   0.49102469913555885   0.025444039112071548   0.8168875466706966   0.8829297825307554   0.2636940404218262   0.703220164181095   0.5097705363625553   0.35112856303434026   0.914749988213113   0.10000184010731242   0.040287724899154824   0.7732779350460826   0.34961098982984173   0.25599815970337036   0.8650327327565148   0.31351396316350094   0.49812821206991753   0.3680182824836477   0.08076759789247288   0.15244813384529374   0.2526762046393169   0.776503037585466   0.3008706866870113   0.3343826925692768   0.761651505503758   0.7510589984733945   0.48398314001631465   0.4514529100385214   0.49795746508193184   0.04783883429229953   0.9742126036537593   0.10032434700418114   0.5832074768688188   0.9478369941849871   0.9339248787546045   0.3270464119580985   0.23359648703897706   0.6918388344816168   0.06889214599808963   0.013532448794597614   0.7354682749690595   0.32382055199796905   0.9881245481056168   0.8610843149493039   0.4827920703297426
0.547317514412503   0.6872538614186054   0.526701622380027   0.7211405648259845   0.7962585159391086   0.20327072140229077   0.07524871234150571   0.22318309974405268   0.7484196816468089   0.2290581177485315   0.9749243653373246   0.6399756228752339   0.8005826874618219   0.295133238993927   0.647877953379226   0.40637913583625684   0.10874385298020514   0.2262410929958374   0.6343455045846285   0.6709108608671973   0.7849233009822361   0.23811654489022066   0.7732611896353245   0.18811879053745473   0.23760578656973308   0.5508626834716153   0.24655956725529746   0.4669782257114702   0.44134727063062457   0.34759196206932447   0.17131085491379175   0.2437951259674175   0.6929275889838156   0.11853384432079296   0.19638648957646718   0.6038195030921837   0.8923449015219936   0.823400605326866   0.5485085361972412   0.1974403672559268   0.7836010485417886   0.5971595123310285   0.9141630316126127   0.5265295063887295   0.9986777475595524   0.3590429674408079   0.14090184197728814   0.33841071585127475   0.7610719609898194   0.8081802839691926   0.8943422747219907   0.8714324901398046   0.3197246903591948   0.4605883218998682   0.723031419808199   0.627637364172387   0.6267971013753793   0.34205447757907526   0.5266449302317318   0.02381786108020342   0.7344521998533856   0.5186538722522093   0.9781363940344907   0.8263774938242766
0.950851151311597   0.9214943599211808   0.06397336242187798   0.29984798743554714   0.9521734037520446   0.5624513924803729   0.9230715204445898   0.9614372715842724   0.1911014427622252   0.7542711085111803   0.028729245722599137   0.09000478144446779   0.8713767524030304   0.29368278661131203   0.3056978259144002   0.46236741727208075   0.24457965102765108   0.9516283090322368   0.7790528956826683   0.4385495561918773   0.5101274511742655   0.4329744367800275   0.8009165016481777   0.6121720623676007   0.5592762998626685   0.5114800768588467   0.7369431392262997   0.31232407493205355   0.6071028961106238   0.9490286843784738   0.8138716187817099   0.3508868033477812   0.4160014533483986   0.19475757586729356   0.7851423730591107   0.26088202190331344   0.5446247009453682   0.9010747892559815   0.4794445471447106   0.7985146046312327   0.30004504991771713   0.9494464802237447   0.7003916514620422   0.35996504843935534   0.7899175987434517   0.5164720434437172   0.8994751498138644   0.7477929860717547   0.23064129888078322   0.004991966584870534   0.16253201058756478   0.4354689111397011   0.6235384027701594   0.05596328220639672   0.3486603918058549   0.08458210779191987   0.2075369494217608   0.8612057063391032   0.5635180187467442   0.8237000858886064   0.6629122484763925   0.9601309170831216   0.08407347160203361   0.02518548125737375
0.36286719855867544   0.010684436859376917   0.3836818201399914   0.6652204328180183   0.5729495998152238   0.49421239341565965   0.48420667032612696   0.9174274467462638   0.3423083009344406   0.48922042683078915   0.3216746597385622   0.48195853560656265   0.7187698981642812   0.4332571446243924   0.9730142679327073   0.3973764278146428   0.5112329487425205   0.5720514382852893   0.40949624918596306   0.5736763419260363   0.8483207002661278   0.6119205212021676   0.32542277758392946   0.5484908606686626   0.48545350170745244   0.6012360843427907   0.941740957443938   0.8832704278506442   0.9125039018922286   0.10702369092713102   0.4575342871178111   0.9658429811043805   0.5701956009577881   0.6178032640963419   0.13585962737924892   0.48388444549781784   0.8514257027935069   0.18454611947194946   0.1628453594465417   0.08650801768317505   0.3401927540509865   0.6124946811866602   0.7533491102605786   0.5128316757571387   0.4918720537848586   0.0005741599844926069   0.42792633267664915   0.9643408150884761   0.006418552077406195   0.39933807564170193   0.4861853752327111   0.08107038723783189   0.09391465018517754   0.2923143847145709   0.028651088114900036   0.11522740613345141   0.5237190492273894   0.674511120618229   0.8927914607356511   0.6313429606356336   0.6722933464338826   0.48996500114627956   0.7299461012891094   0.5448349429524585
0.33210059238289613   0.8774703199596193   0.9765969910285308   0.03200326719531984   0.8402285385980375   0.8768961599751267   0.5486706583518817   0.06766245210684374   0.8338099865206313   0.47755808433342484   0.06248528311917057   0.9865920648690119   0.7398953363354538   0.18524369961885392   0.03383419500427054   0.8713646587355605   0.21617628710806427   0.5107325790006249   0.14104273426861944   0.24002169809992685   0.5438829406741816   0.020767577854345343   0.41109663297951   0.6951867551474683   0.21178234829128556   0.143297257894726   0.4344996419509792   0.6631834879521484   0.3715538096932481   0.26640109791959926   0.8858289835990975   0.5955210358453047   0.5377438231726168   0.7888430135861745   0.8233437004799269   0.608928970976293   0.797848486837163   0.6035993139673206   0.7895095054756563   0.7375643122407325   0.5816721997290988   0.09286673496669563   0.6484667712070369   0.49754261414080564   0.03778925905491711   0.07209915711235029   0.23737013822752695   0.8023558589933373   0.8260069107636315   0.9288018992176242   0.8028704962765478   0.13917237104118882   0.45445310107038345   0.662400801298025   0.9170415126774504   0.543651335195884   0.9167092778977667   0.8735577877118506   0.09369781219752345   0.9347223642195912   0.11886079106060363   0.26995847374453   0.3041883067218671   0.19715805197885872
