3 9
A 1 2 3
B 1 5 7
C 19 20 20
D 1 5 3
E 5 5 2
F 10 8 9
G 2 10 9
H 20 15 19
I 20 2 19
